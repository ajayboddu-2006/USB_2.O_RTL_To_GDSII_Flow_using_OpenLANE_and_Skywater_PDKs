VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO usb
  CLASS BLOCK ;
  FOREIGN usb ;
  ORIGIN 0.000 0.000 ;
  SIZE 177.545 BY 188.265 ;
  PIN clk_48
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END clk_48
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 184.265 149.870 188.265 ;
    END
  END data_in[0]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END data_in[1]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 184.265 80.870 188.265 ;
    END
  END data_in[2]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 184.265 14.170 188.265 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 173.545 166.640 177.545 167.240 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 173.545 105.440 177.545 106.040 ;
    END
  END data_in[7]
  PIN data_in_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 173.545 125.840 177.545 126.440 ;
    END
  END data_in_valid
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 184.265 67.070 188.265 ;
    END
  END data_out[0]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 184.265 53.270 188.265 ;
    END
  END data_out[1]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 184.265 122.270 188.265 ;
    END
  END data_out[2]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END data_out[7]
  PIN data_strobe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END data_strobe
  PIN data_toggle
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 184.265 39.470 188.265 ;
    END
  END data_toggle
  PIN direction_in
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END direction_in
  PIN endpoint[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END endpoint[0]
  PIN endpoint[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 173.545 64.640 177.545 65.240 ;
    END
  END endpoint[1]
  PIN endpoint[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END endpoint[2]
  PIN endpoint[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END endpoint[3]
  PIN handshake[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END handshake[0]
  PIN handshake[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END handshake[1]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 184.265 136.070 188.265 ;
    END
  END rst_n
  PIN rx_j
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 184.265 25.670 188.265 ;
    END
  END rx_j
  PIN rx_se0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 173.545 146.240 177.545 146.840 ;
    END
  END rx_se0
  PIN setup
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 173.545 3.440 177.545 4.040 ;
    END
  END setup
  PIN success
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 184.265 108.470 188.265 ;
    END
  END success
  PIN transaction_active
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END transaction_active
  PIN tx_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 173.545 85.040 177.545 85.640 ;
    END
  END tx_en
  PIN tx_j
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END tx_j
  PIN tx_se0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END tx_se0
  PIN usb_address[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END usb_address[0]
  PIN usb_address[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 184.265 163.670 188.265 ;
    END
  END usb_address[1]
  PIN usb_address[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 184.265 94.670 188.265 ;
    END
  END usb_address[2]
  PIN usb_address[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 173.545 44.240 177.545 44.840 ;
    END
  END usb_address[3]
  PIN usb_address[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END usb_address[4]
  PIN usb_address[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END usb_address[5]
  PIN usb_address[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 184.265 175.170 188.265 ;
    END
  END usb_address[6]
  PIN usb_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 173.545 23.840 177.545 24.440 ;
    END
  END usb_rst
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 143.105 10.640 144.705 177.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 87.750 10.640 89.350 177.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 32.395 10.640 33.995 177.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 148.105 171.580 149.705 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 92.800 171.580 94.400 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 37.495 171.580 39.095 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 115.425 10.640 117.025 177.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 60.075 10.640 61.675 177.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 120.455 171.580 122.055 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 65.145 171.580 66.745 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 171.580 176.885 ;
      LAYER met1 ;
        RECT 2.370 10.640 175.190 177.440 ;
      LAYER met2 ;
        RECT 2.400 183.985 13.610 184.265 ;
        RECT 14.450 183.985 25.110 184.265 ;
        RECT 25.950 183.985 38.910 184.265 ;
        RECT 39.750 183.985 52.710 184.265 ;
        RECT 53.550 183.985 66.510 184.265 ;
        RECT 67.350 183.985 80.310 184.265 ;
        RECT 81.150 183.985 94.110 184.265 ;
        RECT 94.950 183.985 107.910 184.265 ;
        RECT 108.750 183.985 121.710 184.265 ;
        RECT 122.550 183.985 135.510 184.265 ;
        RECT 136.350 183.985 149.310 184.265 ;
        RECT 150.150 183.985 163.110 184.265 ;
        RECT 163.950 183.985 174.610 184.265 ;
        RECT 2.400 4.280 175.160 183.985 ;
        RECT 2.950 3.555 13.610 4.280 ;
        RECT 14.450 3.555 27.410 4.280 ;
        RECT 28.250 3.555 41.210 4.280 ;
        RECT 42.050 3.555 55.010 4.280 ;
        RECT 55.850 3.555 68.810 4.280 ;
        RECT 69.650 3.555 82.610 4.280 ;
        RECT 83.450 3.555 96.410 4.280 ;
        RECT 97.250 3.555 110.210 4.280 ;
        RECT 111.050 3.555 124.010 4.280 ;
        RECT 124.850 3.555 137.810 4.280 ;
        RECT 138.650 3.555 151.610 4.280 ;
        RECT 152.450 3.555 163.110 4.280 ;
        RECT 163.950 3.555 175.160 4.280 ;
      LAYER met3 ;
        RECT 4.400 183.240 173.545 184.105 ;
        RECT 4.000 167.640 173.545 183.240 ;
        RECT 4.000 166.240 173.145 167.640 ;
        RECT 4.000 164.240 173.545 166.240 ;
        RECT 4.400 162.840 173.545 164.240 ;
        RECT 4.000 147.240 173.545 162.840 ;
        RECT 4.000 145.840 173.145 147.240 ;
        RECT 4.000 143.840 173.545 145.840 ;
        RECT 4.400 142.440 173.545 143.840 ;
        RECT 4.000 126.840 173.545 142.440 ;
        RECT 4.000 125.440 173.145 126.840 ;
        RECT 4.000 123.440 173.545 125.440 ;
        RECT 4.400 122.040 173.545 123.440 ;
        RECT 4.000 106.440 173.545 122.040 ;
        RECT 4.000 105.040 173.145 106.440 ;
        RECT 4.000 103.040 173.545 105.040 ;
        RECT 4.400 101.640 173.545 103.040 ;
        RECT 4.000 86.040 173.545 101.640 ;
        RECT 4.000 84.640 173.145 86.040 ;
        RECT 4.000 82.640 173.545 84.640 ;
        RECT 4.400 81.240 173.545 82.640 ;
        RECT 4.000 65.640 173.545 81.240 ;
        RECT 4.000 64.240 173.145 65.640 ;
        RECT 4.000 62.240 173.545 64.240 ;
        RECT 4.400 60.840 173.545 62.240 ;
        RECT 4.000 45.240 173.545 60.840 ;
        RECT 4.000 43.840 173.145 45.240 ;
        RECT 4.000 41.840 173.545 43.840 ;
        RECT 4.400 40.440 173.545 41.840 ;
        RECT 4.000 24.840 173.545 40.440 ;
        RECT 4.000 23.440 173.145 24.840 ;
        RECT 4.000 21.440 173.545 23.440 ;
        RECT 4.400 20.040 173.545 21.440 ;
        RECT 4.000 4.440 173.545 20.040 ;
        RECT 4.000 3.575 173.145 4.440 ;
      LAYER met4 ;
        RECT 62.075 10.640 87.350 177.040 ;
        RECT 89.750 10.640 115.025 177.040 ;
        RECT 117.425 10.640 142.705 177.040 ;
      LAYER met5 ;
        RECT 5.520 96.000 171.580 118.855 ;
        RECT 5.520 68.345 171.580 91.200 ;
        RECT 5.520 40.695 171.580 63.545 ;
  END
END usb
END LIBRARY

