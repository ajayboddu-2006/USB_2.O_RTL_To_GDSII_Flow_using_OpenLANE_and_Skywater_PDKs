magic
tech sky130A
magscale 1 2
timestamp 1738175533
<< checkpaint >>
rect -3932 -3932 39441 41585
<< locali >>
rect 13461 26299 13495 26469
rect 12725 25823 12759 25993
rect 24225 25687 24259 25789
rect 15117 25143 15151 25449
rect 11437 18751 11471 18921
<< viali >>
rect 1593 35241 1627 35275
rect 7205 35241 7239 35275
rect 21741 35241 21775 35275
rect 24501 35241 24535 35275
rect 10609 35173 10643 35207
rect 13369 35173 13403 35207
rect 32597 35173 32631 35207
rect 1409 35105 1443 35139
rect 2789 35105 2823 35139
rect 5089 35105 5123 35139
rect 7389 35105 7423 35139
rect 8217 35105 8251 35139
rect 10793 35105 10827 35139
rect 13553 35105 13587 35139
rect 16313 35105 16347 35139
rect 18889 35105 18923 35139
rect 21833 35105 21867 35139
rect 24593 35105 24627 35139
rect 27353 35105 27387 35139
rect 30021 35105 30055 35139
rect 31953 35105 31987 35139
rect 8033 35037 8067 35071
rect 8125 35037 8159 35071
rect 27169 35037 27203 35071
rect 5273 34969 5307 35003
rect 2973 34901 3007 34935
rect 8585 34901 8619 34935
rect 16129 34901 16163 34935
rect 19073 34901 19107 34935
rect 29837 34901 29871 34935
rect 31769 34901 31803 34935
rect 32505 34901 32539 34935
rect 8401 34697 8435 34731
rect 29377 34697 29411 34731
rect 9827 34629 9861 34663
rect 12081 34629 12115 34663
rect 15209 34629 15243 34663
rect 7757 34561 7791 34595
rect 7941 34561 7975 34595
rect 12633 34561 12667 34595
rect 20867 34561 20901 34595
rect 9689 34493 9723 34527
rect 9965 34493 9999 34527
rect 10149 34493 10183 34527
rect 13829 34493 13863 34527
rect 14085 34493 14119 34527
rect 19073 34493 19107 34527
rect 19441 34493 19475 34527
rect 22661 34493 22695 34527
rect 23029 34493 23063 34527
rect 29469 34493 29503 34527
rect 8033 34357 8067 34391
rect 10149 34357 10183 34391
rect 12449 34357 12483 34391
rect 12541 34357 12575 34391
rect 24455 34357 24489 34391
rect 12265 34153 12299 34187
rect 12633 34153 12667 34187
rect 12725 34153 12759 34187
rect 23305 34153 23339 34187
rect 23765 34153 23799 34187
rect 10140 34085 10174 34119
rect 13461 34017 13495 34051
rect 17141 34017 17175 34051
rect 23673 34017 23707 34051
rect 9873 33949 9907 33983
rect 12817 33949 12851 33983
rect 17509 33949 17543 33983
rect 21005 33949 21039 33983
rect 21373 33949 21407 33983
rect 23949 33949 23983 33983
rect 11253 33813 11287 33847
rect 13553 33813 13587 33847
rect 18935 33813 18969 33847
rect 22799 33813 22833 33847
rect 8217 33609 8251 33643
rect 12817 33609 12851 33643
rect 18153 33609 18187 33643
rect 19441 33609 19475 33643
rect 21649 33609 21683 33643
rect 16129 33541 16163 33575
rect 3893 33473 3927 33507
rect 7665 33473 7699 33507
rect 12173 33473 12207 33507
rect 12357 33473 12391 33507
rect 14381 33473 14415 33507
rect 18797 33473 18831 33507
rect 19901 33473 19935 33507
rect 20085 33473 20119 33507
rect 21005 33473 21039 33507
rect 21189 33473 21223 33507
rect 3709 33405 3743 33439
rect 3801 33405 3835 33439
rect 3985 33405 4019 33439
rect 8677 33405 8711 33439
rect 8953 33405 8987 33439
rect 9505 33405 9539 33439
rect 10517 33405 10551 33439
rect 13277 33405 13311 33439
rect 13461 33405 13495 33439
rect 25329 33405 25363 33439
rect 25697 33405 25731 33439
rect 27905 33405 27939 33439
rect 33609 33405 33643 33439
rect 10333 33337 10367 33371
rect 12449 33337 12483 33371
rect 13369 33337 13403 33371
rect 14657 33337 14691 33371
rect 28181 33337 28215 33371
rect 29929 33337 29963 33371
rect 3525 33269 3559 33303
rect 7757 33269 7791 33303
rect 7849 33269 7883 33303
rect 8769 33269 8803 33303
rect 18521 33269 18555 33303
rect 18613 33269 18647 33303
rect 19809 33269 19843 33303
rect 21281 33269 21315 33303
rect 23903 33269 23937 33303
rect 33425 33269 33459 33303
rect 1593 33065 1627 33099
rect 10517 33065 10551 33099
rect 12449 33065 12483 33099
rect 18199 32997 18233 33031
rect 19993 32997 20027 33031
rect 23581 32997 23615 33031
rect 1409 32929 1443 32963
rect 5650 32929 5684 32963
rect 5917 32929 5951 32963
rect 7685 32929 7719 32963
rect 8401 32929 8435 32963
rect 9597 32929 9631 32963
rect 10057 32929 10091 32963
rect 10517 32929 10551 32963
rect 10701 32929 10735 32963
rect 12817 32929 12851 32963
rect 15117 32929 15151 32963
rect 16405 32929 16439 32963
rect 23434 32929 23468 32963
rect 33425 32929 33459 32963
rect 7941 32861 7975 32895
rect 9873 32861 9907 32895
rect 12909 32861 12943 32895
rect 13001 32861 13035 32895
rect 15209 32861 15243 32895
rect 15301 32861 15335 32895
rect 16773 32861 16807 32895
rect 20140 32861 20174 32895
rect 20361 32861 20395 32895
rect 23213 32861 23247 32895
rect 22937 32793 22971 32827
rect 23305 32793 23339 32827
rect 4537 32725 4571 32759
rect 6561 32725 6595 32759
rect 8493 32725 8527 32759
rect 9735 32725 9769 32759
rect 9965 32725 9999 32759
rect 14749 32725 14783 32759
rect 20269 32725 20303 32759
rect 20453 32725 20487 32759
rect 33517 32725 33551 32759
rect 5089 32521 5123 32555
rect 8309 32521 8343 32555
rect 9045 32521 9079 32555
rect 13093 32521 13127 32555
rect 13553 32521 13587 32555
rect 14841 32521 14875 32555
rect 17969 32453 18003 32487
rect 19349 32453 19383 32487
rect 21603 32453 21637 32487
rect 24777 32453 24811 32487
rect 28917 32453 28951 32487
rect 5733 32385 5767 32419
rect 7481 32385 7515 32419
rect 12541 32385 12575 32419
rect 14013 32385 14047 32419
rect 14105 32385 14139 32419
rect 15301 32385 15335 32419
rect 15393 32385 15427 32419
rect 18613 32385 18647 32419
rect 22753 32385 22787 32419
rect 24225 32385 24259 32419
rect 26525 32385 26559 32419
rect 29469 32385 29503 32419
rect 3626 32317 3660 32351
rect 3893 32317 3927 32351
rect 5457 32317 5491 32351
rect 8493 32317 8527 32351
rect 8585 32317 8619 32351
rect 9045 32317 9079 32351
rect 9229 32317 9263 32351
rect 9781 32317 9815 32351
rect 10048 32317 10082 32351
rect 13921 32317 13955 32351
rect 15209 32317 15243 32351
rect 19165 32317 19199 32351
rect 19349 32317 19383 32351
rect 19809 32317 19843 32351
rect 20177 32317 20211 32351
rect 22937 32317 22971 32351
rect 24317 32317 24351 32351
rect 30113 32317 30147 32351
rect 8309 32249 8343 32283
rect 18429 32249 18463 32283
rect 24409 32249 24443 32283
rect 26341 32249 26375 32283
rect 30389 32249 30423 32283
rect 2513 32181 2547 32215
rect 5549 32181 5583 32215
rect 6929 32181 6963 32215
rect 7297 32181 7331 32215
rect 7389 32181 7423 32215
rect 11161 32181 11195 32215
rect 12633 32181 12667 32215
rect 12725 32181 12759 32215
rect 18337 32181 18371 32215
rect 22845 32181 22879 32215
rect 23305 32181 23339 32215
rect 25881 32181 25915 32215
rect 26249 32181 26283 32215
rect 29285 32181 29319 32215
rect 29377 32181 29411 32215
rect 31861 32181 31895 32215
rect 3341 31977 3375 32011
rect 5733 31977 5767 32011
rect 7849 31977 7883 32011
rect 9597 31977 9631 32011
rect 10241 31977 10275 32011
rect 12449 31977 12483 32011
rect 13001 31977 13035 32011
rect 15485 31977 15519 32011
rect 19993 31977 20027 32011
rect 20361 31977 20395 32011
rect 20453 31977 20487 32011
rect 27307 31977 27341 32011
rect 30481 31977 30515 32011
rect 30849 31977 30883 32011
rect 6736 31909 6770 31943
rect 15025 31909 15059 31943
rect 29101 31909 29135 31943
rect 32137 31909 32171 31943
rect 3157 31841 3191 31875
rect 4537 31841 4571 31875
rect 5365 31841 5399 31875
rect 6469 31841 6503 31875
rect 9689 31841 9723 31875
rect 10149 31841 10183 31875
rect 10333 31841 10367 31875
rect 12357 31841 12391 31875
rect 13001 31841 13035 31875
rect 13185 31841 13219 31875
rect 15117 31841 15151 31875
rect 16221 31841 16255 31875
rect 23121 31841 23155 31875
rect 25881 31841 25915 31875
rect 29009 31841 29043 31875
rect 2973 31773 3007 31807
rect 4353 31773 4387 31807
rect 4721 31773 4755 31807
rect 5273 31773 5307 31807
rect 5457 31773 5491 31807
rect 5549 31773 5583 31807
rect 14841 31773 14875 31807
rect 16589 31773 16623 31807
rect 20637 31773 20671 31807
rect 21695 31773 21729 31807
rect 23489 31773 23523 31807
rect 25513 31773 25547 31807
rect 29285 31773 29319 31807
rect 30941 31773 30975 31807
rect 31125 31773 31159 31807
rect 31769 31705 31803 31739
rect 18015 31637 18049 31671
rect 28641 31637 28675 31671
rect 31677 31637 31711 31671
rect 13921 31433 13955 31467
rect 17509 31433 17543 31467
rect 22661 31433 22695 31467
rect 18981 31365 19015 31399
rect 4077 31297 4111 31331
rect 4261 31297 4295 31331
rect 12541 31297 12575 31331
rect 18153 31297 18187 31331
rect 18852 31297 18886 31331
rect 19073 31297 19107 31331
rect 23581 31297 23615 31331
rect 28089 31297 28123 31331
rect 31401 31297 31435 31331
rect 3985 31229 4019 31263
rect 5641 31229 5675 31263
rect 5917 31229 5951 31263
rect 6837 31229 6871 31263
rect 7021 31229 7055 31263
rect 9505 31229 9539 31263
rect 10149 31229 10183 31263
rect 10333 31229 10367 31263
rect 12633 31229 12667 31263
rect 13737 31229 13771 31263
rect 13921 31229 13955 31263
rect 15761 31229 15795 31263
rect 17969 31229 18003 31263
rect 22845 31229 22879 31263
rect 23949 31229 23983 31263
rect 27813 31229 27847 31263
rect 31217 31229 31251 31263
rect 9260 31161 9294 31195
rect 15494 31161 15528 31195
rect 17877 31161 17911 31195
rect 18705 31161 18739 31195
rect 3617 31093 3651 31127
rect 5825 31093 5859 31127
rect 7205 31093 7239 31127
rect 8125 31093 8159 31127
rect 10149 31093 10183 31127
rect 12725 31093 12759 31127
rect 13093 31093 13127 31127
rect 14381 31093 14415 31127
rect 19349 31093 19383 31127
rect 25375 31093 25409 31127
rect 29561 31093 29595 31127
rect 30849 31093 30883 31127
rect 31309 31093 31343 31127
rect 6653 30889 6687 30923
rect 11621 30889 11655 30923
rect 12449 30889 12483 30923
rect 14841 30889 14875 30923
rect 17923 30889 17957 30923
rect 23029 30889 23063 30923
rect 23581 30889 23615 30923
rect 24041 30889 24075 30923
rect 32505 30889 32539 30923
rect 12817 30821 12851 30855
rect 31033 30821 31067 30855
rect 3157 30753 3191 30787
rect 5273 30753 5307 30787
rect 5641 30753 5675 30787
rect 5917 30753 5951 30787
rect 6929 30753 6963 30787
rect 7113 30753 7147 30787
rect 10497 30753 10531 30787
rect 12909 30753 12943 30787
rect 14749 30753 14783 30787
rect 20545 30753 20579 30787
rect 22845 30753 22879 30787
rect 23949 30753 23983 30787
rect 27721 30753 27755 30787
rect 30757 30753 30791 30787
rect 2973 30685 3007 30719
rect 3065 30685 3099 30719
rect 3249 30685 3283 30719
rect 4997 30685 5031 30719
rect 6837 30685 6871 30719
rect 7021 30685 7055 30719
rect 10241 30685 10275 30719
rect 13093 30685 13127 30719
rect 16129 30685 16163 30719
rect 16497 30685 16531 30719
rect 20637 30685 20671 30719
rect 20729 30685 20763 30719
rect 24133 30685 24167 30719
rect 25927 30685 25961 30719
rect 27353 30685 27387 30719
rect 2789 30549 2823 30583
rect 20177 30549 20211 30583
rect 4813 30345 4847 30379
rect 10057 30345 10091 30379
rect 24455 30345 24489 30379
rect 6837 30277 6871 30311
rect 13185 30277 13219 30311
rect 13737 30277 13771 30311
rect 15117 30277 15151 30311
rect 18245 30277 18279 30311
rect 26065 30277 26099 30311
rect 7481 30209 7515 30243
rect 14289 30209 14323 30243
rect 15209 30209 15243 30243
rect 18705 30209 18739 30243
rect 18889 30209 18923 30243
rect 21097 30209 21131 30243
rect 22661 30209 22695 30243
rect 23029 30209 23063 30243
rect 26617 30209 26651 30243
rect 29377 30209 29411 30243
rect 1409 30141 1443 30175
rect 1676 30141 1710 30175
rect 3709 30141 3743 30175
rect 4169 30141 4203 30175
rect 4537 30141 4571 30175
rect 7205 30141 7239 30175
rect 8769 30141 8803 30175
rect 9965 30141 9999 30175
rect 10149 30141 10183 30175
rect 10609 30141 10643 30175
rect 10793 30141 10827 30175
rect 11437 30141 11471 30175
rect 13093 30141 13127 30175
rect 13277 30141 13311 30175
rect 14197 30141 14231 30175
rect 14933 30141 14967 30175
rect 15025 30141 15059 30175
rect 18613 30141 18647 30175
rect 21465 30141 21499 30175
rect 25329 30141 25363 30175
rect 26525 30141 26559 30175
rect 29193 30141 29227 30175
rect 29837 30141 29871 30175
rect 30021 30141 30055 30175
rect 7297 30073 7331 30107
rect 10701 30073 10735 30107
rect 14105 30073 14139 30107
rect 2789 30005 2823 30039
rect 8861 30005 8895 30039
rect 11253 30005 11287 30039
rect 19671 30005 19705 30039
rect 25513 30005 25547 30039
rect 26433 30005 26467 30039
rect 2973 29801 3007 29835
rect 5641 29801 5675 29835
rect 9781 29801 9815 29835
rect 10977 29801 11011 29835
rect 12633 29801 12667 29835
rect 14933 29801 14967 29835
rect 4721 29733 4755 29767
rect 11345 29733 11379 29767
rect 12541 29733 12575 29767
rect 16414 29733 16448 29767
rect 3157 29665 3191 29699
rect 4629 29665 4663 29699
rect 5733 29665 5767 29699
rect 5917 29665 5951 29699
rect 7757 29665 7791 29699
rect 9505 29665 9539 29699
rect 10241 29665 10275 29699
rect 10425 29665 10459 29699
rect 14749 29665 14783 29699
rect 25237 29665 25271 29699
rect 26065 29665 26099 29699
rect 26157 29665 26191 29699
rect 26249 29665 26283 29699
rect 27997 29665 28031 29699
rect 28365 29665 28399 29699
rect 28825 29665 28859 29699
rect 3341 29597 3375 29631
rect 4905 29597 4939 29631
rect 7481 29597 7515 29631
rect 7665 29597 7699 29631
rect 9781 29597 9815 29631
rect 10333 29597 10367 29631
rect 11437 29597 11471 29631
rect 11621 29597 11655 29631
rect 12817 29597 12851 29631
rect 16681 29597 16715 29631
rect 17233 29597 17267 29631
rect 17601 29597 17635 29631
rect 19027 29597 19061 29631
rect 21097 29597 21131 29631
rect 21465 29597 21499 29631
rect 30665 29597 30699 29631
rect 30941 29597 30975 29631
rect 9597 29529 9631 29563
rect 12173 29529 12207 29563
rect 25881 29529 25915 29563
rect 27905 29529 27939 29563
rect 4261 29461 4295 29495
rect 8125 29461 8159 29495
rect 15301 29461 15335 29495
rect 22891 29461 22925 29495
rect 25329 29461 25363 29495
rect 32413 29461 32447 29495
rect 1961 29257 1995 29291
rect 8033 29257 8067 29291
rect 9873 29257 9907 29291
rect 12449 29257 12483 29291
rect 12725 29257 12759 29291
rect 18337 29257 18371 29291
rect 23397 29257 23431 29291
rect 25329 29257 25363 29291
rect 25513 29257 25547 29291
rect 30665 29257 30699 29291
rect 5549 29189 5583 29223
rect 8493 29189 8527 29223
rect 26525 29189 26559 29223
rect 33425 29189 33459 29223
rect 3249 29121 3283 29155
rect 3433 29121 3467 29155
rect 7389 29121 7423 29155
rect 7573 29121 7607 29155
rect 8953 29121 8987 29155
rect 9137 29121 9171 29155
rect 13277 29121 13311 29155
rect 14381 29121 14415 29155
rect 18797 29121 18831 29155
rect 18981 29121 19015 29155
rect 27997 29121 28031 29155
rect 31217 29121 31251 29155
rect 1777 29053 1811 29087
rect 3341 29053 3375 29087
rect 3525 29053 3559 29087
rect 4077 29053 4111 29087
rect 4261 29053 4295 29087
rect 4353 29053 4387 29087
rect 5273 29053 5307 29087
rect 5365 29053 5399 29087
rect 5641 29053 5675 29087
rect 7665 29053 7699 29087
rect 9781 29053 9815 29087
rect 10517 29053 10551 29087
rect 10701 29053 10735 29087
rect 12633 29053 12667 29087
rect 13093 29053 13127 29087
rect 17325 29053 17359 29087
rect 17509 29053 17543 29087
rect 18705 29053 18739 29087
rect 20361 29053 20395 29087
rect 20545 29053 20579 29087
rect 23581 29053 23615 29087
rect 24225 29053 24259 29087
rect 24409 29053 24443 29087
rect 26341 29053 26375 29087
rect 31033 29053 31067 29087
rect 33609 29053 33643 29087
rect 13185 28985 13219 29019
rect 17693 28985 17727 29019
rect 25145 28985 25179 29019
rect 28273 28985 28307 29019
rect 31125 28985 31159 29019
rect 3065 28917 3099 28951
rect 5089 28917 5123 28951
rect 8861 28917 8895 28951
rect 10609 28917 10643 28951
rect 14565 28917 14599 28951
rect 14657 28917 14691 28951
rect 15025 28917 15059 28951
rect 20361 28917 20395 28951
rect 24317 28917 24351 28951
rect 25350 28917 25384 28951
rect 29745 28917 29779 28951
rect 3157 28713 3191 28747
rect 6193 28713 6227 28747
rect 8585 28713 8619 28747
rect 9781 28713 9815 28747
rect 10241 28713 10275 28747
rect 12357 28713 12391 28747
rect 14749 28713 14783 28747
rect 19073 28713 19107 28747
rect 21189 28713 21223 28747
rect 23673 28713 23707 28747
rect 25442 28713 25476 28747
rect 26111 28713 26145 28747
rect 28825 28713 28859 28747
rect 30665 28713 30699 28747
rect 2044 28645 2078 28679
rect 5080 28645 5114 28679
rect 7021 28645 7055 28679
rect 15117 28645 15151 28679
rect 19993 28645 20027 28679
rect 20177 28645 20211 28679
rect 22109 28645 22143 28679
rect 25237 28645 25271 28679
rect 29193 28645 29227 28679
rect 32404 28645 32438 28679
rect 1777 28577 1811 28611
rect 4813 28577 4847 28611
rect 8401 28577 8435 28611
rect 8585 28577 8619 28611
rect 9873 28577 9907 28611
rect 10977 28577 11011 28611
rect 11233 28577 11267 28611
rect 12817 28577 12851 28611
rect 13001 28577 13035 28611
rect 13645 28577 13679 28611
rect 16773 28577 16807 28611
rect 19073 28577 19107 28611
rect 20269 28577 20303 28611
rect 20913 28577 20947 28611
rect 21005 28577 21039 28611
rect 21281 28577 21315 28611
rect 22017 28577 22051 28611
rect 22201 28577 22235 28611
rect 23949 28577 23983 28611
rect 24133 28577 24167 28611
rect 27905 28577 27939 28611
rect 31033 28577 31067 28611
rect 7113 28509 7147 28543
rect 7297 28509 7331 28543
rect 9597 28509 9631 28543
rect 13737 28509 13771 28543
rect 15209 28509 15243 28543
rect 15301 28509 15335 28543
rect 16589 28509 16623 28543
rect 18797 28509 18831 28543
rect 21097 28509 21131 28543
rect 23857 28509 23891 28543
rect 24041 28509 24075 28543
rect 27537 28509 27571 28543
rect 29285 28509 29319 28543
rect 29469 28509 29503 28543
rect 30481 28509 30515 28543
rect 30941 28509 30975 28543
rect 32137 28509 32171 28543
rect 18981 28441 19015 28475
rect 6653 28373 6687 28407
rect 12909 28373 12943 28407
rect 16957 28373 16991 28407
rect 20085 28373 20119 28407
rect 25421 28373 25455 28407
rect 25605 28373 25639 28407
rect 33517 28373 33551 28407
rect 3709 28169 3743 28203
rect 4445 28169 4479 28203
rect 5549 28169 5583 28203
rect 11069 28169 11103 28203
rect 13001 28169 13035 28203
rect 20269 28169 20303 28203
rect 25789 28169 25823 28203
rect 30205 28169 30239 28203
rect 31677 28169 31711 28203
rect 17417 28101 17451 28135
rect 20913 28101 20947 28135
rect 24961 28101 24995 28135
rect 25559 28101 25593 28135
rect 25697 28101 25731 28135
rect 9873 28033 9907 28067
rect 14749 28033 14783 28067
rect 17785 28033 17819 28067
rect 19165 28033 19199 28067
rect 21557 28033 21591 28067
rect 26433 28033 26467 28067
rect 28457 28033 28491 28067
rect 5365 27965 5399 27999
rect 8125 27965 8159 27999
rect 8309 27965 8343 27999
rect 10057 27965 10091 27999
rect 10241 27965 10275 27999
rect 10977 27965 11011 27999
rect 11161 27965 11195 27999
rect 12817 27965 12851 27999
rect 13001 27965 13035 27999
rect 14657 27965 14691 27999
rect 18889 27965 18923 27999
rect 20177 27965 20211 27999
rect 20361 27965 20395 27999
rect 20821 27965 20855 27999
rect 21005 27965 21039 27999
rect 21465 27965 21499 27999
rect 23949 27965 23983 27999
rect 24225 27965 24259 27999
rect 24685 27965 24719 27999
rect 24777 27965 24811 27999
rect 24961 27965 24995 27999
rect 25421 27965 25455 27999
rect 25881 27965 25915 27999
rect 26341 27965 26375 27999
rect 26525 27965 26559 27999
rect 30849 27965 30883 27999
rect 31033 27965 31067 27999
rect 31493 27965 31527 27999
rect 3617 27897 3651 27931
rect 4353 27897 4387 27931
rect 5181 27897 5215 27931
rect 17969 27897 18003 27931
rect 23029 27897 23063 27931
rect 24133 27897 24167 27931
rect 28733 27897 28767 27931
rect 8217 27829 8251 27863
rect 14197 27829 14231 27863
rect 14565 27829 14599 27863
rect 17877 27829 17911 27863
rect 18521 27829 18555 27863
rect 18981 27829 19015 27863
rect 23121 27829 23155 27863
rect 23765 27829 23799 27863
rect 30665 27829 30699 27863
rect 4721 27625 4755 27659
rect 13093 27625 13127 27659
rect 14749 27625 14783 27659
rect 15117 27625 15151 27659
rect 21005 27625 21039 27659
rect 25237 27625 25271 27659
rect 28825 27625 28859 27659
rect 32576 27625 32610 27659
rect 10057 27557 10091 27591
rect 10425 27557 10459 27591
rect 11437 27557 11471 27591
rect 13553 27557 13587 27591
rect 20729 27557 20763 27591
rect 21649 27557 21683 27591
rect 31708 27557 31742 27591
rect 32781 27557 32815 27591
rect 2973 27489 3007 27523
rect 4629 27489 4663 27523
rect 7225 27489 7259 27523
rect 8217 27489 8251 27523
rect 8401 27489 8435 27523
rect 8493 27489 8527 27523
rect 10241 27489 10275 27523
rect 11345 27489 11379 27523
rect 11529 27489 11563 27523
rect 11989 27489 12023 27523
rect 12173 27489 12207 27523
rect 13461 27489 13495 27523
rect 17233 27489 17267 27523
rect 19993 27489 20027 27523
rect 20913 27489 20947 27523
rect 21005 27489 21039 27523
rect 21833 27489 21867 27523
rect 21923 27489 21957 27523
rect 22385 27489 22419 27523
rect 22477 27489 22511 27523
rect 22661 27489 22695 27523
rect 24409 27489 24443 27523
rect 25237 27489 25271 27523
rect 25421 27489 25455 27523
rect 29009 27489 29043 27523
rect 29285 27489 29319 27523
rect 2881 27421 2915 27455
rect 3065 27421 3099 27455
rect 3157 27421 3191 27455
rect 4905 27421 4939 27455
rect 7481 27421 7515 27455
rect 13645 27421 13679 27455
rect 15209 27421 15243 27455
rect 15301 27421 15335 27455
rect 17601 27421 17635 27455
rect 31953 27421 31987 27455
rect 4261 27353 4295 27387
rect 6101 27353 6135 27387
rect 8217 27353 8251 27387
rect 24593 27353 24627 27387
rect 29101 27353 29135 27387
rect 29193 27353 29227 27387
rect 2697 27285 2731 27319
rect 12081 27285 12115 27319
rect 19027 27285 19061 27319
rect 20177 27285 20211 27319
rect 21925 27285 21959 27319
rect 22845 27285 22879 27319
rect 30573 27285 30607 27319
rect 32413 27285 32447 27319
rect 32597 27285 32631 27319
rect 10425 27081 10459 27115
rect 12357 27081 12391 27115
rect 13461 27081 13495 27115
rect 14657 27081 14691 27115
rect 24777 27081 24811 27115
rect 13369 27013 13403 27047
rect 14105 27013 14139 27047
rect 16405 27013 16439 27047
rect 17601 27013 17635 27047
rect 24225 27013 24259 27047
rect 1501 26945 1535 26979
rect 3985 26945 4019 26979
rect 7941 26945 7975 26979
rect 8125 26945 8159 26979
rect 13553 26945 13587 26979
rect 18153 26945 18187 26979
rect 19441 26945 19475 26979
rect 20913 26945 20947 26979
rect 21097 26945 21131 26979
rect 22753 26945 22787 26979
rect 27905 26945 27939 26979
rect 29837 26945 29871 26979
rect 30757 26945 30791 26979
rect 1768 26877 1802 26911
rect 4537 26877 4571 26911
rect 7849 26877 7883 26911
rect 8677 26877 8711 26911
rect 8953 26877 8987 26911
rect 9505 26877 9539 26911
rect 10609 26877 10643 26911
rect 10885 26877 10919 26911
rect 12449 26877 12483 26911
rect 12909 26877 12943 26911
rect 13277 26877 13311 26911
rect 14013 26877 14047 26911
rect 14841 26877 14875 26911
rect 15025 26877 15059 26911
rect 15292 26877 15326 26911
rect 17325 26877 17359 26911
rect 17877 26877 17911 26911
rect 18981 26877 19015 26911
rect 20821 26877 20855 26911
rect 22569 26877 22603 26911
rect 22661 26877 22695 26911
rect 22937 26877 22971 26911
rect 23397 26877 23431 26911
rect 23581 26877 23615 26911
rect 24041 26877 24075 26911
rect 24317 26877 24351 26911
rect 24593 26877 24627 26911
rect 27997 26877 28031 26911
rect 30113 26877 30147 26911
rect 31024 26877 31058 26911
rect 33149 26877 33183 26911
rect 33333 26877 33367 26911
rect 3801 26809 3835 26843
rect 4804 26809 4838 26843
rect 10793 26809 10827 26843
rect 23489 26809 23523 26843
rect 33057 26809 33091 26843
rect 2881 26741 2915 26775
rect 3341 26741 3375 26775
rect 3709 26741 3743 26775
rect 5917 26741 5951 26775
rect 7481 26741 7515 26775
rect 8769 26741 8803 26775
rect 13093 26741 13127 26775
rect 20453 26741 20487 26775
rect 22845 26741 22879 26775
rect 24409 26741 24443 26775
rect 28365 26741 28399 26775
rect 32137 26741 32171 26775
rect 2973 26537 3007 26571
rect 4905 26537 4939 26571
rect 7481 26537 7515 26571
rect 8401 26537 8435 26571
rect 10057 26537 10091 26571
rect 16773 26537 16807 26571
rect 19073 26537 19107 26571
rect 27813 26537 27847 26571
rect 33149 26537 33183 26571
rect 7389 26469 7423 26503
rect 11345 26469 11379 26503
rect 12265 26469 12299 26503
rect 12470 26469 12504 26503
rect 13461 26469 13495 26503
rect 13553 26469 13587 26503
rect 14749 26469 14783 26503
rect 16681 26469 16715 26503
rect 22523 26469 22557 26503
rect 26341 26469 26375 26503
rect 3157 26401 3191 26435
rect 5089 26401 5123 26435
rect 5181 26401 5215 26435
rect 8309 26401 8343 26435
rect 10425 26401 10459 26435
rect 11621 26401 11655 26435
rect 3341 26333 3375 26367
rect 5549 26333 5583 26367
rect 7205 26333 7239 26367
rect 10517 26333 10551 26367
rect 10701 26333 10735 26367
rect 11253 26333 11287 26367
rect 11805 26333 11839 26367
rect 13737 26401 13771 26435
rect 14933 26401 14967 26435
rect 15577 26401 15611 26435
rect 16957 26401 16991 26435
rect 18705 26401 18739 26435
rect 18889 26401 18923 26435
rect 21097 26401 21131 26435
rect 23121 26401 23155 26435
rect 23305 26401 23339 26435
rect 24133 26401 24167 26435
rect 24317 26401 24351 26435
rect 25329 26401 25363 26435
rect 25513 26401 25547 26435
rect 29377 26401 29411 26435
rect 29561 26401 29595 26435
rect 30941 26401 30975 26435
rect 31309 26401 31343 26435
rect 32036 26401 32070 26435
rect 20729 26333 20763 26367
rect 23029 26333 23063 26367
rect 23949 26333 23983 26367
rect 26065 26333 26099 26367
rect 30757 26333 30791 26367
rect 31769 26333 31803 26367
rect 13461 26265 13495 26299
rect 17141 26265 17175 26299
rect 25513 26265 25547 26299
rect 31217 26265 31251 26299
rect 7849 26197 7883 26231
rect 12449 26197 12483 26231
rect 12633 26197 12667 26231
rect 29469 26197 29503 26231
rect 4905 25993 4939 26027
rect 7941 25993 7975 26027
rect 10517 25993 10551 26027
rect 12725 25993 12759 26027
rect 14565 25993 14599 26027
rect 21051 25993 21085 26027
rect 22845 25993 22879 26027
rect 10977 25925 11011 25959
rect 12173 25925 12207 25959
rect 3433 25857 3467 25891
rect 7297 25857 7331 25891
rect 7481 25857 7515 25891
rect 8953 25857 8987 25891
rect 30941 25925 30975 25959
rect 19625 25857 19659 25891
rect 26341 25857 26375 25891
rect 26525 25857 26559 25891
rect 30205 25857 30239 25891
rect 32045 25857 32079 25891
rect 33333 25857 33367 25891
rect 5089 25789 5123 25823
rect 5365 25789 5399 25823
rect 7573 25789 7607 25823
rect 10333 25789 10367 25823
rect 10517 25789 10551 25823
rect 11161 25789 11195 25823
rect 12081 25789 12115 25823
rect 12265 25789 12299 25823
rect 12725 25789 12759 25823
rect 12817 25789 12851 25823
rect 15209 25789 15243 25823
rect 16129 25789 16163 25823
rect 17325 25789 17359 25823
rect 17509 25789 17543 25823
rect 19257 25789 19291 25823
rect 23029 25789 23063 25823
rect 23305 25789 23339 25823
rect 24225 25789 24259 25823
rect 24317 25789 24351 25823
rect 24593 25789 24627 25823
rect 25329 25789 25363 25823
rect 26249 25789 26283 25823
rect 28181 25789 28215 25823
rect 30757 25789 30791 25823
rect 31401 25789 31435 25823
rect 33057 25789 33091 25823
rect 33241 25789 33275 25823
rect 3157 25721 3191 25755
rect 9137 25721 9171 25755
rect 13093 25721 13127 25755
rect 24685 25721 24719 25755
rect 28457 25721 28491 25755
rect 5273 25653 5307 25687
rect 9045 25653 9079 25687
rect 9505 25653 9539 25687
rect 15209 25653 15243 25687
rect 16037 25653 16071 25687
rect 17417 25653 17451 25687
rect 23213 25653 23247 25687
rect 24225 25653 24259 25687
rect 25237 25653 25271 25687
rect 25881 25653 25915 25687
rect 8125 25449 8159 25483
rect 13093 25449 13127 25483
rect 15117 25449 15151 25483
rect 25421 25449 25455 25483
rect 28549 25449 28583 25483
rect 29469 25449 29503 25483
rect 5043 25381 5077 25415
rect 9689 25381 9723 25415
rect 12817 25381 12851 25415
rect 1777 25313 1811 25347
rect 1961 25313 1995 25347
rect 2513 25313 2547 25347
rect 2605 25313 2639 25347
rect 4721 25313 4755 25347
rect 4813 25313 4847 25347
rect 4905 25313 4939 25347
rect 7389 25313 7423 25347
rect 7941 25313 7975 25347
rect 9873 25313 9907 25347
rect 10885 25313 10919 25347
rect 11161 25313 11195 25347
rect 11253 25313 11287 25347
rect 12449 25313 12483 25347
rect 12541 25313 12575 25347
rect 12725 25313 12759 25347
rect 12909 25313 12943 25347
rect 1869 25245 1903 25279
rect 2697 25245 2731 25279
rect 2789 25245 2823 25279
rect 5181 25245 5215 25279
rect 7113 25245 7147 25279
rect 10609 25177 10643 25211
rect 23949 25381 23983 25415
rect 26534 25381 26568 25415
rect 32965 25381 32999 25415
rect 15476 25313 15510 25347
rect 18714 25313 18748 25347
rect 23213 25313 23247 25347
rect 23489 25313 23523 25347
rect 24133 25313 24167 25347
rect 24317 25313 24351 25347
rect 28181 25313 28215 25347
rect 28335 25313 28369 25347
rect 29377 25313 29411 25347
rect 29561 25313 29595 25347
rect 30941 25313 30975 25347
rect 31585 25313 31619 25347
rect 31769 25313 31803 25347
rect 32229 25313 32263 25347
rect 33517 25313 33551 25347
rect 15209 25245 15243 25279
rect 18981 25245 19015 25279
rect 26801 25245 26835 25279
rect 32321 25177 32355 25211
rect 2973 25109 3007 25143
rect 4537 25109 4571 25143
rect 5641 25109 5675 25143
rect 9505 25109 9539 25143
rect 15117 25109 15151 25143
rect 16589 25109 16623 25143
rect 17601 25109 17635 25143
rect 23397 25109 23431 25143
rect 5181 24905 5215 24939
rect 6837 24905 6871 24939
rect 8309 24905 8343 24939
rect 16221 24905 16255 24939
rect 30757 24905 30791 24939
rect 7297 24769 7331 24803
rect 7481 24769 7515 24803
rect 9413 24769 9447 24803
rect 10793 24769 10827 24803
rect 12081 24769 12115 24803
rect 15577 24769 15611 24803
rect 16313 24769 16347 24803
rect 18889 24769 18923 24803
rect 23489 24769 23523 24803
rect 33333 24769 33367 24803
rect 2789 24701 2823 24735
rect 4454 24701 4488 24735
rect 4721 24701 4755 24735
rect 5181 24701 5215 24735
rect 5365 24701 5399 24735
rect 7205 24701 7239 24735
rect 8309 24701 8343 24735
rect 9229 24701 9263 24735
rect 10241 24701 10275 24735
rect 10701 24701 10735 24735
rect 10885 24701 10919 24735
rect 12265 24701 12299 24735
rect 12357 24701 12391 24735
rect 13645 24701 13679 24735
rect 15301 24701 15335 24735
rect 16037 24701 16071 24735
rect 16129 24701 16163 24735
rect 17509 24701 17543 24735
rect 17785 24701 17819 24735
rect 17969 24701 18003 24735
rect 21281 24701 21315 24735
rect 21557 24701 21591 24735
rect 22661 24701 22695 24735
rect 23581 24701 23615 24735
rect 23765 24701 23799 24735
rect 24133 24701 24167 24735
rect 25053 24701 25087 24735
rect 27997 24701 28031 24735
rect 28273 24701 28307 24735
rect 29745 24701 29779 24735
rect 29929 24701 29963 24735
rect 30297 24701 30331 24735
rect 32137 24701 32171 24735
rect 33057 24701 33091 24735
rect 33241 24701 33275 24735
rect 2544 24633 2578 24667
rect 9321 24633 9355 24667
rect 14841 24633 14875 24667
rect 15393 24633 15427 24667
rect 19165 24633 19199 24667
rect 21465 24633 21499 24667
rect 31892 24633 31926 24667
rect 1409 24565 1443 24599
rect 3341 24565 3375 24599
rect 8861 24565 8895 24599
rect 10149 24565 10183 24599
rect 12081 24565 12115 24599
rect 13829 24565 13863 24599
rect 17325 24565 17359 24599
rect 20637 24565 20671 24599
rect 21373 24565 21407 24599
rect 22753 24565 22787 24599
rect 25237 24565 25271 24599
rect 28095 24565 28129 24599
rect 28181 24565 28215 24599
rect 29929 24565 29963 24599
rect 1593 24361 1627 24395
rect 13001 24361 13035 24395
rect 18153 24361 18187 24395
rect 18705 24361 18739 24395
rect 20177 24361 20211 24395
rect 23510 24361 23544 24395
rect 24317 24361 24351 24395
rect 29193 24361 29227 24395
rect 31217 24361 31251 24395
rect 2789 24293 2823 24327
rect 6285 24293 6319 24327
rect 8217 24293 8251 24327
rect 11253 24293 11287 24327
rect 18857 24293 18891 24327
rect 19073 24293 19107 24327
rect 23305 24293 23339 24327
rect 27169 24293 27203 24327
rect 1409 24225 1443 24259
rect 2145 24225 2179 24259
rect 3157 24225 3191 24259
rect 3341 24225 3375 24259
rect 4445 24225 4479 24259
rect 5181 24225 5215 24259
rect 6193 24225 6227 24259
rect 8033 24225 8067 24259
rect 12173 24225 12207 24259
rect 12909 24225 12943 24259
rect 16404 24225 16438 24259
rect 16497 24225 16531 24259
rect 17141 24225 17175 24259
rect 17969 24225 18003 24259
rect 18153 24225 18187 24259
rect 19993 24225 20027 24259
rect 24133 24225 24167 24259
rect 24317 24225 24351 24259
rect 25513 24225 25547 24259
rect 25881 24225 25915 24259
rect 25973 24225 26007 24259
rect 29101 24225 29135 24259
rect 29285 24225 29319 24259
rect 31309 24225 31343 24259
rect 5273 24157 5307 24191
rect 11529 24157 11563 24191
rect 12449 24157 12483 24191
rect 17233 24157 17267 24191
rect 21005 24157 21039 24191
rect 21373 24157 21407 24191
rect 26893 24157 26927 24191
rect 28641 24157 28675 24191
rect 31217 24157 31251 24191
rect 31861 24157 31895 24191
rect 32137 24157 32171 24191
rect 3157 24089 3191 24123
rect 4629 24089 4663 24123
rect 8401 24089 8435 24123
rect 16129 24089 16163 24123
rect 17509 24089 17543 24123
rect 2237 24021 2271 24055
rect 9781 24021 9815 24055
rect 12265 24021 12299 24055
rect 12357 24021 12391 24055
rect 18889 24021 18923 24055
rect 22799 24021 22833 24055
rect 23489 24021 23523 24055
rect 23673 24021 23707 24055
rect 25329 24021 25363 24055
rect 30757 24021 30791 24055
rect 33609 24021 33643 24055
rect 2697 23817 2731 23851
rect 9229 23817 9263 23851
rect 10517 23817 10551 23851
rect 12357 23817 12391 23851
rect 19441 23817 19475 23851
rect 25329 23817 25363 23851
rect 3525 23749 3559 23783
rect 9873 23749 9907 23783
rect 29469 23749 29503 23783
rect 4445 23681 4479 23715
rect 4997 23681 5031 23715
rect 8033 23681 8067 23715
rect 8217 23681 8251 23715
rect 8769 23681 8803 23715
rect 13461 23681 13495 23715
rect 30849 23681 30883 23715
rect 2789 23613 2823 23647
rect 4813 23613 4847 23647
rect 5365 23613 5399 23647
rect 5825 23613 5859 23647
rect 8309 23613 8343 23647
rect 8953 23613 8987 23647
rect 9045 23613 9079 23647
rect 9321 23613 9355 23647
rect 9781 23613 9815 23647
rect 9965 23613 9999 23647
rect 10425 23613 10459 23647
rect 10609 23613 10643 23647
rect 12173 23613 12207 23647
rect 12265 23613 12299 23647
rect 13185 23613 13219 23647
rect 19717 23613 19751 23647
rect 22937 23613 22971 23647
rect 23397 23613 23431 23647
rect 23857 23613 23891 23647
rect 24225 23613 24259 23647
rect 25145 23613 25179 23647
rect 25421 23613 25455 23647
rect 28365 23613 28399 23647
rect 28549 23613 28583 23647
rect 29653 23613 29687 23647
rect 30481 23613 30515 23647
rect 31585 23613 31619 23647
rect 31861 23613 31895 23647
rect 3341 23545 3375 23579
rect 12449 23545 12483 23579
rect 19441 23545 19475 23579
rect 24317 23545 24351 23579
rect 25666 23545 25700 23579
rect 31401 23545 31435 23579
rect 8033 23477 8067 23511
rect 14933 23477 14967 23511
rect 19625 23477 19659 23511
rect 22753 23477 22787 23511
rect 26801 23477 26835 23511
rect 28181 23477 28215 23511
rect 31769 23477 31803 23511
rect 11989 23273 12023 23307
rect 14841 23273 14875 23307
rect 17233 23273 17267 23307
rect 17877 23273 17911 23307
rect 20913 23273 20947 23307
rect 25329 23273 25363 23307
rect 28733 23273 28767 23307
rect 32873 23273 32907 23307
rect 33241 23273 33275 23307
rect 10149 23205 10183 23239
rect 12081 23205 12115 23239
rect 16120 23205 16154 23239
rect 18981 23205 19015 23239
rect 20545 23205 20579 23239
rect 23549 23205 23583 23239
rect 23765 23205 23799 23239
rect 25789 23205 25823 23239
rect 5089 23137 5123 23171
rect 5917 23137 5951 23171
rect 7113 23137 7147 23171
rect 7665 23137 7699 23171
rect 10057 23137 10091 23171
rect 10333 23137 10367 23171
rect 10609 23137 10643 23171
rect 10793 23137 10827 23171
rect 11897 23137 11931 23171
rect 12173 23137 12207 23171
rect 12633 23137 12667 23171
rect 12817 23137 12851 23171
rect 14933 23137 14967 23171
rect 15853 23137 15887 23171
rect 17693 23137 17727 23171
rect 18797 23137 18831 23171
rect 19073 23137 19107 23171
rect 20361 23137 20395 23171
rect 20637 23137 20671 23171
rect 20729 23137 20763 23171
rect 22385 23137 22419 23171
rect 25697 23137 25731 23171
rect 27813 23137 27847 23171
rect 30665 23137 30699 23171
rect 1409 23069 1443 23103
rect 1685 23069 1719 23103
rect 5365 23069 5399 23103
rect 5641 23069 5675 23103
rect 21741 23069 21775 23103
rect 25881 23069 25915 23103
rect 28825 23069 28859 23103
rect 28917 23069 28951 23103
rect 30941 23069 30975 23103
rect 32413 23069 32447 23103
rect 33333 23069 33367 23103
rect 33425 23069 33459 23103
rect 4813 23001 4847 23035
rect 8033 23001 8067 23035
rect 3157 22933 3191 22967
rect 12725 22933 12759 22967
rect 18797 22933 18831 22967
rect 23397 22933 23431 22967
rect 23581 22933 23615 22967
rect 27629 22933 27663 22967
rect 28365 22933 28399 22967
rect 3433 22729 3467 22763
rect 4169 22729 4203 22763
rect 6929 22729 6963 22763
rect 10977 22729 11011 22763
rect 13001 22729 13035 22763
rect 15853 22729 15887 22763
rect 19533 22729 19567 22763
rect 26801 22729 26835 22763
rect 30021 22729 30055 22763
rect 30849 22729 30883 22763
rect 5825 22661 5859 22695
rect 13093 22661 13127 22695
rect 23765 22661 23799 22695
rect 4813 22593 4847 22627
rect 8401 22593 8435 22627
rect 8677 22593 8711 22627
rect 13185 22593 13219 22627
rect 14105 22593 14139 22627
rect 18797 22593 18831 22627
rect 19717 22593 19751 22627
rect 20545 22593 20579 22627
rect 24685 22593 24719 22627
rect 28549 22593 28583 22627
rect 31401 22593 31435 22627
rect 2697 22525 2731 22559
rect 2881 22525 2915 22559
rect 3341 22525 3375 22559
rect 3525 22525 3559 22559
rect 4353 22525 4387 22559
rect 4445 22525 4479 22559
rect 5549 22525 5583 22559
rect 5825 22525 5859 22559
rect 9137 22525 9171 22559
rect 11069 22525 11103 22559
rect 12081 22525 12115 22559
rect 12265 22525 12299 22559
rect 12909 22525 12943 22559
rect 19073 22525 19107 22559
rect 19533 22525 19567 22559
rect 19901 22525 19935 22559
rect 20361 22525 20395 22559
rect 20729 22525 20763 22559
rect 22753 22525 22787 22559
rect 22937 22525 22971 22559
rect 23397 22525 23431 22559
rect 23489 22525 23523 22559
rect 23857 22525 23891 22559
rect 23949 22525 23983 22559
rect 24409 22525 24443 22559
rect 26709 22525 26743 22559
rect 28273 22525 28307 22559
rect 31309 22525 31343 22559
rect 4721 22457 4755 22491
rect 14381 22457 14415 22491
rect 22845 22457 22879 22491
rect 2789 22389 2823 22423
rect 9321 22389 9355 22423
rect 12173 22389 12207 22423
rect 17325 22389 17359 22423
rect 19809 22389 19843 22423
rect 20453 22389 20487 22423
rect 20637 22389 20671 22423
rect 26157 22389 26191 22423
rect 31217 22389 31251 22423
rect 4813 22185 4847 22219
rect 10977 22185 11011 22219
rect 12357 22185 12391 22219
rect 16681 22117 16715 22151
rect 22373 22117 22407 22151
rect 30665 22117 30699 22151
rect 30870 22117 30904 22151
rect 2973 22049 3007 22083
rect 4721 22049 4755 22083
rect 4905 22049 4939 22083
rect 5365 22049 5399 22083
rect 5549 22049 5583 22083
rect 6469 22049 6503 22083
rect 6929 22049 6963 22083
rect 7205 22049 7239 22083
rect 11161 22049 11195 22083
rect 12357 22049 12391 22083
rect 13369 22049 13403 22083
rect 16405 22049 16439 22083
rect 16589 22049 16623 22083
rect 22753 22049 22787 22083
rect 23397 22049 23431 22083
rect 25973 22049 26007 22083
rect 26433 22049 26467 22083
rect 27077 22049 27111 22083
rect 27445 22049 27479 22083
rect 27721 22049 27755 22083
rect 28273 22049 28307 22083
rect 28641 22049 28675 22083
rect 29285 22049 29319 22083
rect 31677 22049 31711 22083
rect 32045 22049 32079 22083
rect 32689 22049 32723 22083
rect 2697 21981 2731 22015
rect 7113 21981 7147 22015
rect 11989 21981 12023 22015
rect 12541 21981 12575 22015
rect 13645 21981 13679 22015
rect 20177 21981 20211 22015
rect 20453 21981 20487 22015
rect 23765 21981 23799 22015
rect 26709 21981 26743 22015
rect 31493 21981 31527 22015
rect 13461 21913 13495 21947
rect 31033 21913 31067 21947
rect 2789 21845 2823 21879
rect 2881 21845 2915 21879
rect 5549 21845 5583 21879
rect 13553 21845 13587 21879
rect 21925 21845 21959 21879
rect 28365 21845 28399 21879
rect 30849 21845 30883 21879
rect 11161 21641 11195 21675
rect 12817 21641 12851 21675
rect 19993 21641 20027 21675
rect 21281 21641 21315 21675
rect 21649 21641 21683 21675
rect 23213 21641 23247 21675
rect 24409 21641 24443 21675
rect 25329 21641 25363 21675
rect 25513 21641 25547 21675
rect 24777 21573 24811 21607
rect 28457 21573 28491 21607
rect 30573 21573 30607 21607
rect 1685 21505 1719 21539
rect 3157 21505 3191 21539
rect 4813 21505 4847 21539
rect 4997 21505 5031 21539
rect 8861 21505 8895 21539
rect 14381 21505 14415 21539
rect 17785 21505 17819 21539
rect 22569 21505 22603 21539
rect 31493 21505 31527 21539
rect 31677 21505 31711 21539
rect 1409 21437 1443 21471
rect 3893 21437 3927 21471
rect 4077 21437 4111 21471
rect 8033 21437 8067 21471
rect 8493 21437 8527 21471
rect 8677 21437 8711 21471
rect 9413 21437 9447 21471
rect 12081 21437 12115 21471
rect 12269 21437 12303 21471
rect 12360 21437 12394 21471
rect 12449 21437 12483 21471
rect 12633 21437 12667 21471
rect 13829 21437 13863 21471
rect 14473 21437 14507 21471
rect 14565 21437 14599 21471
rect 15025 21437 15059 21471
rect 15485 21437 15519 21471
rect 17969 21437 18003 21471
rect 20085 21437 20119 21471
rect 21465 21437 21499 21471
rect 21649 21437 21683 21471
rect 22937 21437 22971 21471
rect 23029 21437 23063 21471
rect 24593 21437 24627 21471
rect 24869 21437 24903 21471
rect 27997 21437 28031 21471
rect 28273 21437 28307 21471
rect 30389 21437 30423 21471
rect 33609 21437 33643 21471
rect 9689 21369 9723 21403
rect 22707 21369 22741 21403
rect 22845 21369 22879 21403
rect 25697 21369 25731 21403
rect 29193 21369 29227 21403
rect 31769 21369 31803 21403
rect 3985 21301 4019 21335
rect 5089 21301 5123 21335
rect 5457 21301 5491 21335
rect 18153 21301 18187 21335
rect 25492 21301 25526 21335
rect 29101 21301 29135 21335
rect 32137 21301 32171 21335
rect 33425 21301 33459 21335
rect 4997 21097 5031 21131
rect 7297 21097 7331 21131
rect 11437 21097 11471 21131
rect 15853 21097 15887 21131
rect 17693 21097 17727 21131
rect 2973 21029 3007 21063
rect 6469 21029 6503 21063
rect 8217 21029 8251 21063
rect 8309 21029 8343 21063
rect 9505 21029 9539 21063
rect 9689 21029 9723 21063
rect 11989 21029 12023 21063
rect 22477 21029 22511 21063
rect 24041 21029 24075 21063
rect 25789 21029 25823 21063
rect 32137 21029 32171 21063
rect 3157 20961 3191 20995
rect 3249 20961 3283 20995
rect 4261 20961 4295 20995
rect 5181 20961 5215 20995
rect 5365 20961 5399 20995
rect 5733 20961 5767 20995
rect 6377 20961 6411 20995
rect 7205 20961 7239 20995
rect 8125 20961 8159 20995
rect 8447 20961 8481 20995
rect 10333 20961 10367 20995
rect 10517 20961 10551 20995
rect 11253 20961 11287 20995
rect 11437 20961 11471 20995
rect 11897 20961 11931 20995
rect 12357 20961 12391 20995
rect 12725 20961 12759 20995
rect 15025 20961 15059 20995
rect 16580 20961 16614 20995
rect 18705 20961 18739 20995
rect 20361 20961 20395 20995
rect 22385 20961 22419 20995
rect 22569 20961 22603 20995
rect 23305 20961 23339 20995
rect 23489 20961 23523 20995
rect 23949 20961 23983 20995
rect 25605 20961 25639 20995
rect 26525 20961 26559 20995
rect 27261 20961 27295 20995
rect 29110 20961 29144 20995
rect 30849 20961 30883 20995
rect 4905 20893 4939 20927
rect 5641 20893 5675 20927
rect 8585 20893 8619 20927
rect 12449 20893 12483 20927
rect 12633 20893 12667 20927
rect 14933 20893 14967 20927
rect 16313 20893 16347 20927
rect 18981 20893 19015 20927
rect 20269 20893 20303 20927
rect 25421 20893 25455 20927
rect 29377 20893 29411 20927
rect 30941 20893 30975 20927
rect 31125 20893 31159 20927
rect 31861 20893 31895 20927
rect 33609 20893 33643 20927
rect 2973 20825 3007 20859
rect 4353 20825 4387 20859
rect 10333 20825 10367 20859
rect 18889 20825 18923 20859
rect 27077 20825 27111 20859
rect 7941 20757 7975 20791
rect 9873 20757 9907 20791
rect 18521 20757 18555 20791
rect 19993 20757 20027 20791
rect 20177 20757 20211 20791
rect 23305 20757 23339 20791
rect 26433 20757 26467 20791
rect 27997 20757 28031 20791
rect 30481 20757 30515 20791
rect 2973 20553 3007 20587
rect 3341 20553 3375 20587
rect 3985 20553 4019 20587
rect 6929 20553 6963 20587
rect 10517 20553 10551 20587
rect 10977 20553 11011 20587
rect 12265 20553 12299 20587
rect 19441 20553 19475 20587
rect 25973 20553 26007 20587
rect 26617 20553 26651 20587
rect 28089 20553 28123 20587
rect 31309 20553 31343 20587
rect 32137 20553 32171 20587
rect 17417 20485 17451 20519
rect 1777 20417 1811 20451
rect 3433 20417 3467 20451
rect 8401 20417 8435 20451
rect 8677 20417 8711 20451
rect 18061 20417 18095 20451
rect 28641 20417 28675 20451
rect 29837 20417 29871 20451
rect 3157 20349 3191 20383
rect 3893 20349 3927 20383
rect 5089 20349 5123 20383
rect 5549 20349 5583 20383
rect 5733 20349 5767 20383
rect 9597 20349 9631 20383
rect 10517 20349 10551 20383
rect 10701 20349 10735 20383
rect 10793 20349 10827 20383
rect 11069 20349 11103 20383
rect 12173 20349 12207 20383
rect 12357 20349 12391 20383
rect 13369 20349 13403 20383
rect 13553 20349 13587 20383
rect 14013 20349 14047 20383
rect 14197 20349 14231 20383
rect 17325 20349 17359 20383
rect 17509 20349 17543 20383
rect 18328 20349 18362 20383
rect 20729 20349 20763 20383
rect 21281 20349 21315 20383
rect 23029 20349 23063 20383
rect 23489 20349 23523 20383
rect 23765 20349 23799 20383
rect 24685 20349 24719 20383
rect 25053 20349 25087 20383
rect 25145 20349 25179 20383
rect 25605 20349 25639 20383
rect 25789 20349 25823 20383
rect 26433 20349 26467 20383
rect 28457 20349 28491 20383
rect 29561 20349 29595 20383
rect 31769 20349 31803 20383
rect 31953 20349 31987 20383
rect 1961 20281 1995 20315
rect 5641 20281 5675 20315
rect 9689 20281 9723 20315
rect 15853 20281 15887 20315
rect 16037 20281 16071 20315
rect 22845 20281 22879 20315
rect 24777 20281 24811 20315
rect 24869 20281 24903 20315
rect 4997 20213 5031 20247
rect 13461 20213 13495 20247
rect 14105 20213 14139 20247
rect 20177 20213 20211 20247
rect 24501 20213 24535 20247
rect 28549 20213 28583 20247
rect 4926 20009 4960 20043
rect 5089 20009 5123 20043
rect 5825 20009 5859 20043
rect 6837 20009 6871 20043
rect 16497 20009 16531 20043
rect 17785 20009 17819 20043
rect 26525 20009 26559 20043
rect 2973 19941 3007 19975
rect 4721 19941 4755 19975
rect 12541 19941 12575 19975
rect 24225 19941 24259 19975
rect 27077 19941 27111 19975
rect 2513 19873 2547 19907
rect 3157 19873 3191 19907
rect 3341 19873 3375 19907
rect 6009 19873 6043 19907
rect 6745 19873 6779 19907
rect 9781 19873 9815 19907
rect 10149 19873 10183 19907
rect 10517 19873 10551 19907
rect 10701 19873 10735 19907
rect 11253 19873 11287 19907
rect 12173 19873 12207 19907
rect 12357 19873 12391 19907
rect 13001 19873 13035 19907
rect 14749 19873 14783 19907
rect 14933 19873 14967 19907
rect 15025 19873 15059 19907
rect 15163 19873 15197 19907
rect 16037 19873 16071 19907
rect 16773 19873 16807 19907
rect 16865 19873 16899 19907
rect 16957 19873 16991 19907
rect 17141 19873 17175 19907
rect 17601 19873 17635 19907
rect 17877 19873 17911 19907
rect 22753 19873 22787 19907
rect 22937 19873 22971 19907
rect 24317 19873 24351 19907
rect 25237 19873 25271 19907
rect 25375 19873 25409 19907
rect 25605 19873 25639 19907
rect 26433 19873 26467 19907
rect 27261 19873 27295 19907
rect 27445 19873 27479 19907
rect 28549 19873 28583 19907
rect 2237 19805 2271 19839
rect 10241 19805 10275 19839
rect 20361 19805 20395 19839
rect 20637 19805 20671 19839
rect 28273 19805 28307 19839
rect 28457 19805 28491 19839
rect 31861 19805 31895 19839
rect 32137 19805 32171 19839
rect 13185 19737 13219 19771
rect 2329 19669 2363 19703
rect 2421 19669 2455 19703
rect 4905 19669 4939 19703
rect 15393 19669 15427 19703
rect 15945 19669 15979 19703
rect 17601 19669 17635 19703
rect 22109 19669 22143 19703
rect 22753 19669 22787 19703
rect 28917 19669 28951 19703
rect 33609 19669 33643 19703
rect 3157 19465 3191 19499
rect 3985 19465 4019 19499
rect 4537 19465 4571 19499
rect 12265 19465 12299 19499
rect 13185 19465 13219 19499
rect 13553 19465 13587 19499
rect 17785 19465 17819 19499
rect 25053 19465 25087 19499
rect 9965 19397 9999 19431
rect 14933 19397 14967 19431
rect 15071 19397 15105 19431
rect 33149 19397 33183 19431
rect 1685 19329 1719 19363
rect 5641 19329 5675 19363
rect 7113 19329 7147 19363
rect 14841 19329 14875 19363
rect 15393 19329 15427 19363
rect 16405 19329 16439 19363
rect 20729 19329 20763 19363
rect 20913 19329 20947 19363
rect 22845 19329 22879 19363
rect 23581 19329 23615 19363
rect 31033 19329 31067 19363
rect 31217 19329 31251 19363
rect 33517 19329 33551 19363
rect 1409 19261 1443 19295
rect 4537 19261 4571 19295
rect 4721 19261 4755 19295
rect 4813 19261 4847 19295
rect 5273 19261 5307 19295
rect 5549 19261 5583 19295
rect 6837 19261 6871 19295
rect 9045 19261 9079 19295
rect 9229 19261 9263 19295
rect 9597 19261 9631 19295
rect 9781 19261 9815 19295
rect 10057 19261 10091 19295
rect 10517 19261 10551 19295
rect 10609 19261 10643 19295
rect 12173 19261 12207 19295
rect 12449 19261 12483 19295
rect 13369 19261 13403 19295
rect 13553 19261 13587 19295
rect 15485 19261 15519 19295
rect 15853 19261 15887 19295
rect 16129 19261 16163 19295
rect 16313 19261 16347 19295
rect 19901 19261 19935 19295
rect 20177 19261 20211 19295
rect 21005 19261 21039 19295
rect 21557 19261 21591 19295
rect 21649 19261 21683 19295
rect 22661 19261 22695 19295
rect 23305 19261 23339 19295
rect 25605 19261 25639 19295
rect 26525 19261 26559 19295
rect 26617 19261 26651 19295
rect 26801 19261 26835 19295
rect 29570 19261 29604 19295
rect 29837 19261 29871 19295
rect 3709 19193 3743 19227
rect 14473 19193 14507 19227
rect 15209 19193 15243 19227
rect 15301 19193 15335 19227
rect 15577 19193 15611 19227
rect 15669 19193 15703 19227
rect 18061 19193 18095 19227
rect 20729 19193 20763 19227
rect 30941 19193 30975 19227
rect 8585 19125 8619 19159
rect 15945 19125 15979 19159
rect 20085 19125 20119 19159
rect 25697 19125 25731 19159
rect 26525 19125 26559 19159
rect 28457 19125 28491 19159
rect 30573 19125 30607 19159
rect 33057 19125 33091 19159
rect 2421 18921 2455 18955
rect 4721 18921 4755 18955
rect 5641 18921 5675 18955
rect 9781 18921 9815 18955
rect 11437 18921 11471 18955
rect 32689 18921 32723 18955
rect 33057 18921 33091 18955
rect 4873 18853 4907 18887
rect 5089 18853 5123 18887
rect 8401 18853 8435 18887
rect 2421 18785 2455 18819
rect 2605 18785 2639 18819
rect 3341 18785 3375 18819
rect 5549 18785 5583 18819
rect 5733 18785 5767 18819
rect 8309 18785 8343 18819
rect 8493 18785 8527 18819
rect 9689 18785 9723 18819
rect 9873 18785 9907 18819
rect 10793 18785 10827 18819
rect 13461 18853 13495 18887
rect 16775 18853 16809 18887
rect 26801 18853 26835 18887
rect 28733 18853 28767 18887
rect 30757 18853 30791 18887
rect 11529 18785 11563 18819
rect 13645 18785 13679 18819
rect 13829 18785 13863 18819
rect 15025 18785 15059 18819
rect 15761 18785 15795 18819
rect 15945 18785 15979 18819
rect 18797 18785 18831 18819
rect 19165 18785 19199 18819
rect 19901 18785 19935 18819
rect 20085 18785 20119 18819
rect 20177 18785 20211 18819
rect 25237 18785 25271 18819
rect 25973 18785 26007 18819
rect 26157 18785 26191 18819
rect 26709 18785 26743 18819
rect 26985 18785 27019 18819
rect 28181 18785 28215 18819
rect 28365 18785 28399 18819
rect 30481 18785 30515 18819
rect 10517 18717 10551 18751
rect 11437 18717 11471 18751
rect 12357 18717 12391 18751
rect 12449 18717 12483 18751
rect 12725 18717 12759 18751
rect 12909 18717 12943 18751
rect 15209 18717 15243 18751
rect 18981 18717 19015 18751
rect 19625 18717 19659 18751
rect 19809 18717 19843 18751
rect 20361 18717 20395 18751
rect 25513 18717 25547 18751
rect 26065 18717 26099 18751
rect 32229 18717 32263 18751
rect 33149 18717 33183 18751
rect 33241 18717 33275 18751
rect 18797 18649 18831 18683
rect 25329 18649 25363 18683
rect 27905 18649 27939 18683
rect 3157 18581 3191 18615
rect 4905 18581 4939 18615
rect 10609 18581 10643 18615
rect 10701 18581 10735 18615
rect 11621 18581 11655 18615
rect 18061 18581 18095 18615
rect 19717 18581 19751 18615
rect 25421 18581 25455 18615
rect 27169 18581 27203 18615
rect 27997 18581 28031 18615
rect 4077 18377 4111 18411
rect 10885 18377 10919 18411
rect 16313 18377 16347 18411
rect 17601 18377 17635 18411
rect 22661 18377 22695 18411
rect 26249 18377 26283 18411
rect 27813 18377 27847 18411
rect 30573 18377 30607 18411
rect 14841 18241 14875 18275
rect 19073 18241 19107 18275
rect 19349 18241 19383 18275
rect 21649 18241 21683 18275
rect 24409 18241 24443 18275
rect 24869 18241 24903 18275
rect 2513 18173 2547 18207
rect 2697 18173 2731 18207
rect 2973 18173 3007 18207
rect 4905 18173 4939 18207
rect 4997 18173 5031 18207
rect 5181 18173 5215 18207
rect 5273 18173 5307 18207
rect 7113 18173 7147 18207
rect 7665 18173 7699 18207
rect 9137 18173 9171 18207
rect 9229 18173 9263 18207
rect 9439 18173 9473 18207
rect 9597 18173 9631 18207
rect 10241 18173 10275 18207
rect 10333 18173 10367 18207
rect 11161 18173 11195 18207
rect 12357 18173 12391 18207
rect 12449 18173 12483 18207
rect 12817 18173 12851 18207
rect 13277 18173 13311 18207
rect 13737 18173 13771 18207
rect 15025 18173 15059 18207
rect 15393 18173 15427 18207
rect 16405 18173 16439 18207
rect 25136 18173 25170 18207
rect 27905 18173 27939 18207
rect 28089 18173 28123 18207
rect 28641 18173 28675 18207
rect 30389 18173 30423 18207
rect 3065 18105 3099 18139
rect 4056 18105 4090 18139
rect 4261 18105 4295 18139
rect 6929 18105 6963 18139
rect 9321 18105 9355 18139
rect 10885 18105 10919 18139
rect 12081 18105 12115 18139
rect 21373 18105 21407 18139
rect 24133 18105 24167 18139
rect 3893 18037 3927 18071
rect 4721 18037 4755 18071
rect 8953 18037 8987 18071
rect 11069 18037 11103 18071
rect 19901 18037 19935 18071
rect 1869 17833 1903 17867
rect 2973 17833 3007 17867
rect 17877 17833 17911 17867
rect 20821 17833 20855 17867
rect 22201 17833 22235 17867
rect 26617 17833 26651 17867
rect 3065 17765 3099 17799
rect 12909 17765 12943 17799
rect 15853 17765 15887 17799
rect 1777 17697 1811 17731
rect 1961 17697 1995 17731
rect 4353 17697 4387 17731
rect 4537 17697 4571 17731
rect 4997 17697 5031 17731
rect 5457 17697 5491 17731
rect 5917 17697 5951 17731
rect 6193 17697 6227 17731
rect 6377 17697 6411 17731
rect 7481 17697 7515 17731
rect 10425 17697 10459 17731
rect 12817 17697 12851 17731
rect 13001 17697 13035 17731
rect 14749 17697 14783 17731
rect 14841 17697 14875 17731
rect 15117 17697 15151 17731
rect 17785 17697 17819 17731
rect 20545 17697 20579 17731
rect 21281 17697 21315 17731
rect 21465 17697 21499 17731
rect 21925 17697 21959 17731
rect 22661 17697 22695 17731
rect 22845 17697 22879 17731
rect 26525 17697 26559 17731
rect 26709 17697 26743 17731
rect 27353 17697 27387 17731
rect 27997 17697 28031 17731
rect 31861 17697 31895 17731
rect 2881 17629 2915 17663
rect 4445 17629 4479 17663
rect 10057 17629 10091 17663
rect 12541 17629 12575 17663
rect 12633 17629 12667 17663
rect 15577 17629 15611 17663
rect 20821 17629 20855 17663
rect 21373 17629 21407 17663
rect 22201 17629 22235 17663
rect 22753 17629 22787 17663
rect 27261 17629 27295 17663
rect 27813 17629 27847 17663
rect 28273 17629 28307 17663
rect 32137 17629 32171 17663
rect 6469 17561 6503 17595
rect 2513 17493 2547 17527
rect 7389 17493 7423 17527
rect 11851 17493 11885 17527
rect 13277 17493 13311 17527
rect 17325 17493 17359 17527
rect 20637 17493 20671 17527
rect 22017 17493 22051 17527
rect 33609 17493 33643 17527
rect 2789 17289 2823 17323
rect 4721 17289 4755 17323
rect 4905 17289 4939 17323
rect 5733 17289 5767 17323
rect 9965 17289 9999 17323
rect 11161 17289 11195 17323
rect 28089 17289 28123 17323
rect 7389 17153 7423 17187
rect 8493 17153 8527 17187
rect 10793 17153 10827 17187
rect 14749 17153 14783 17187
rect 15117 17153 15151 17187
rect 15209 17153 15243 17187
rect 21649 17153 21683 17187
rect 25605 17153 25639 17187
rect 26065 17153 26099 17187
rect 30573 17153 30607 17187
rect 31401 17153 31435 17187
rect 2513 17085 2547 17119
rect 2605 17085 2639 17119
rect 5181 17085 5215 17119
rect 5641 17085 5675 17119
rect 5825 17085 5859 17119
rect 7205 17085 7239 17119
rect 8217 17085 8251 17119
rect 10977 17085 11011 17119
rect 12541 17085 12575 17119
rect 13093 17085 13127 17119
rect 13461 17085 13495 17119
rect 13645 17085 13679 17119
rect 14013 17085 14047 17119
rect 14933 17085 14967 17119
rect 15025 17085 15059 17119
rect 19257 17085 19291 17119
rect 19717 17085 19751 17119
rect 19901 17085 19935 17119
rect 21465 17085 21499 17119
rect 24961 17085 24995 17119
rect 25697 17085 25731 17119
rect 26525 17085 26559 17119
rect 26709 17085 26743 17119
rect 27997 17085 28031 17119
rect 28181 17085 28215 17119
rect 28825 17085 28859 17119
rect 31217 17085 31251 17119
rect 31861 17085 31895 17119
rect 32045 17085 32079 17119
rect 33425 17085 33459 17119
rect 12449 17017 12483 17051
rect 15761 17017 15795 17051
rect 16129 17017 16163 17051
rect 18981 17017 19015 17051
rect 24685 17017 24719 17051
rect 25973 17017 26007 17051
rect 29101 17017 29135 17051
rect 33609 17017 33643 17051
rect 6837 16949 6871 16983
rect 7297 16949 7331 16983
rect 17509 16949 17543 16983
rect 19809 16949 19843 16983
rect 23213 16949 23247 16983
rect 25421 16949 25455 16983
rect 26525 16949 26559 16983
rect 31033 16949 31067 16983
rect 31953 16949 31987 16983
rect 5549 16745 5583 16779
rect 7941 16745 7975 16779
rect 11897 16745 11931 16779
rect 12541 16745 12575 16779
rect 14841 16745 14875 16779
rect 15761 16745 15795 16779
rect 20545 16745 20579 16779
rect 32045 16745 32079 16779
rect 3065 16677 3099 16711
rect 6828 16677 6862 16711
rect 18245 16677 18279 16711
rect 21097 16677 21131 16711
rect 26985 16677 27019 16711
rect 30849 16677 30883 16711
rect 2968 16609 3002 16643
rect 3157 16609 3191 16643
rect 3341 16609 3375 16643
rect 5641 16609 5675 16643
rect 11805 16609 11839 16643
rect 12449 16609 12483 16643
rect 12633 16609 12667 16643
rect 13461 16609 13495 16643
rect 13737 16609 13771 16643
rect 14749 16609 14783 16643
rect 14933 16609 14967 16643
rect 15761 16609 15795 16643
rect 15945 16609 15979 16643
rect 16405 16609 16439 16643
rect 16589 16609 16623 16643
rect 17233 16609 17267 16643
rect 19073 16609 19107 16643
rect 20269 16609 20303 16643
rect 21005 16609 21039 16643
rect 21189 16609 21223 16643
rect 25237 16609 25271 16643
rect 25421 16609 25455 16643
rect 25973 16609 26007 16643
rect 26157 16609 26191 16643
rect 26709 16609 26743 16643
rect 30573 16609 30607 16643
rect 30757 16609 30791 16643
rect 31401 16609 31435 16643
rect 31585 16609 31619 16643
rect 31677 16609 31711 16643
rect 31769 16609 31803 16643
rect 32505 16609 32539 16643
rect 32686 16609 32720 16643
rect 32781 16609 32815 16643
rect 33425 16609 33459 16643
rect 33517 16609 33551 16643
rect 6561 16541 6595 16575
rect 20545 16541 20579 16575
rect 25329 16541 25363 16575
rect 26985 16541 27019 16575
rect 13553 16473 13587 16507
rect 26801 16473 26835 16507
rect 3341 16405 3375 16439
rect 16405 16405 16439 16439
rect 17141 16405 17175 16439
rect 20361 16405 20395 16439
rect 26157 16405 26191 16439
rect 4813 16201 4847 16235
rect 14105 16201 14139 16235
rect 15209 16201 15243 16235
rect 18797 16201 18831 16235
rect 19533 16201 19567 16235
rect 22661 16201 22695 16235
rect 26249 16201 26283 16235
rect 27905 16201 27939 16235
rect 30113 16201 30147 16235
rect 11161 16133 11195 16167
rect 18889 16133 18923 16167
rect 3433 16065 3467 16099
rect 9689 16065 9723 16099
rect 18705 16065 18739 16099
rect 21005 16065 21039 16099
rect 21281 16065 21315 16099
rect 22845 16065 22879 16099
rect 23397 16065 23431 16099
rect 1409 15997 1443 16031
rect 4169 15997 4203 16031
rect 4445 15997 4479 16031
rect 5181 15997 5215 16031
rect 7297 15997 7331 16031
rect 9873 15997 9907 16031
rect 10885 15997 10919 16031
rect 10977 15997 11011 16031
rect 12449 15997 12483 16031
rect 12909 15997 12943 16031
rect 13921 15997 13955 16031
rect 14197 15997 14231 16031
rect 16037 15997 16071 16031
rect 18981 15997 19015 16031
rect 22569 15997 22603 16031
rect 23305 15997 23339 16031
rect 23489 15997 23523 16031
rect 25513 15997 25547 16031
rect 25697 15997 25731 16031
rect 26157 15997 26191 16031
rect 26341 15997 26375 16031
rect 29018 15997 29052 16031
rect 29285 15997 29319 16031
rect 30389 15997 30423 16031
rect 30478 15997 30512 16031
rect 30573 15997 30607 16031
rect 30757 15997 30791 16031
rect 31769 15997 31803 16031
rect 33609 15997 33643 16031
rect 1685 15929 1719 15963
rect 7573 15929 7607 15963
rect 11161 15929 11195 15963
rect 15025 15929 15059 15963
rect 15241 15929 15275 15963
rect 25329 15929 25363 15963
rect 31953 15929 31987 15963
rect 33517 15929 33551 15963
rect 9045 15861 9079 15895
rect 10057 15861 10091 15895
rect 12265 15861 12299 15895
rect 13001 15861 13035 15895
rect 15393 15861 15427 15895
rect 15945 15861 15979 15895
rect 22845 15861 22879 15895
rect 32137 15861 32171 15895
rect 2881 15657 2915 15691
rect 16405 15657 16439 15691
rect 23489 15657 23523 15691
rect 33609 15657 33643 15691
rect 8493 15589 8527 15623
rect 9689 15589 9723 15623
rect 10425 15589 10459 15623
rect 17325 15589 17359 15623
rect 22017 15589 22051 15623
rect 31217 15589 31251 15623
rect 31401 15589 31435 15623
rect 32137 15589 32171 15623
rect 3065 15521 3099 15555
rect 3341 15521 3375 15555
rect 7665 15521 7699 15555
rect 11069 15521 11103 15555
rect 11161 15521 11195 15555
rect 11437 15521 11471 15555
rect 12817 15521 12851 15555
rect 13645 15521 13679 15555
rect 15393 15521 15427 15555
rect 15577 15521 15611 15555
rect 16221 15521 16255 15555
rect 17095 15521 17129 15555
rect 17233 15521 17267 15555
rect 17417 15521 17451 15555
rect 21741 15521 21775 15555
rect 23949 15521 23983 15555
rect 25513 15521 25547 15555
rect 25973 15521 26007 15555
rect 26157 15521 26191 15555
rect 26801 15521 26835 15555
rect 26985 15521 27019 15555
rect 27885 15521 27919 15555
rect 3249 15453 3283 15487
rect 6377 15453 6411 15487
rect 6653 15453 6687 15487
rect 7849 15453 7883 15487
rect 11345 15453 11379 15487
rect 12541 15453 12575 15487
rect 12633 15453 12667 15487
rect 12725 15453 12759 15487
rect 15301 15453 15335 15487
rect 16957 15453 16991 15487
rect 25237 15453 25271 15487
rect 27629 15453 27663 15487
rect 31861 15453 31895 15487
rect 8309 15385 8343 15419
rect 12357 15385 12391 15419
rect 4905 15317 4939 15351
rect 7481 15317 7515 15351
rect 10885 15317 10919 15351
rect 13461 15317 13495 15351
rect 15761 15317 15795 15351
rect 17601 15317 17635 15351
rect 24041 15317 24075 15351
rect 25329 15317 25363 15351
rect 25421 15317 25455 15351
rect 26065 15317 26099 15351
rect 26893 15317 26927 15351
rect 29009 15317 29043 15351
rect 31033 15317 31067 15351
rect 31217 15317 31251 15351
rect 12173 15113 12207 15147
rect 13185 15113 13219 15147
rect 25605 15113 25639 15147
rect 26617 15113 26651 15147
rect 26709 15113 26743 15147
rect 30757 15113 30791 15147
rect 31861 15113 31895 15147
rect 20729 15045 20763 15079
rect 1685 14977 1719 15011
rect 3985 14977 4019 15011
rect 4077 14977 4111 15011
rect 4721 14977 4755 15011
rect 5457 14977 5491 15011
rect 10517 14977 10551 15011
rect 10793 14977 10827 15011
rect 14565 14977 14599 15011
rect 17601 14977 17635 15011
rect 20913 14977 20947 15011
rect 24225 14977 24259 15011
rect 26801 14977 26835 15011
rect 29009 14977 29043 15011
rect 1409 14909 1443 14943
rect 3893 14909 3927 14943
rect 4353 14909 4387 14943
rect 5549 14909 5583 14943
rect 7849 14909 7883 14943
rect 8217 14909 8251 14943
rect 12265 14909 12299 14943
rect 13093 14909 13127 14943
rect 13461 14909 13495 14943
rect 13737 14909 13771 14943
rect 14197 14909 14231 14943
rect 14381 14909 14415 14943
rect 15485 14909 15519 14943
rect 15761 14909 15795 14943
rect 17325 14909 17359 14943
rect 20637 14909 20671 14943
rect 21557 14909 21591 14943
rect 24492 14909 24526 14943
rect 26525 14909 26559 14943
rect 31217 14909 31251 14943
rect 31401 14909 31435 14943
rect 32137 14909 32171 14943
rect 3433 14841 3467 14875
rect 15853 14841 15887 14875
rect 29285 14841 29319 14875
rect 31309 14841 31343 14875
rect 31861 14841 31895 14875
rect 5181 14773 5215 14807
rect 7297 14773 7331 14807
rect 9045 14773 9079 14807
rect 19073 14773 19107 14807
rect 20913 14773 20947 14807
rect 21465 14773 21499 14807
rect 32045 14773 32079 14807
rect 3157 14569 3191 14603
rect 4261 14569 4295 14603
rect 5181 14569 5215 14603
rect 7389 14569 7423 14603
rect 11161 14569 11195 14603
rect 16037 14569 16071 14603
rect 21741 14569 21775 14603
rect 22293 14569 22327 14603
rect 25329 14569 25363 14603
rect 28089 14569 28123 14603
rect 30849 14569 30883 14603
rect 3341 14501 3375 14535
rect 4424 14501 4458 14535
rect 4629 14501 4663 14535
rect 5368 14501 5402 14535
rect 12449 14501 12483 14535
rect 20269 14501 20303 14535
rect 23029 14501 23063 14535
rect 26249 14501 26283 14535
rect 26954 14501 26988 14535
rect 3065 14433 3099 14467
rect 5089 14433 5123 14467
rect 7297 14433 7331 14467
rect 7481 14433 7515 14467
rect 11069 14433 11103 14467
rect 11345 14433 11379 14467
rect 12357 14433 12391 14467
rect 13369 14433 13403 14467
rect 15209 14433 15243 14467
rect 15393 14433 15427 14467
rect 15945 14433 15979 14467
rect 16589 14433 16623 14467
rect 16773 14433 16807 14467
rect 16957 14433 16991 14467
rect 18061 14433 18095 14467
rect 18797 14433 18831 14467
rect 18981 14433 19015 14467
rect 19993 14433 20027 14467
rect 22201 14433 22235 14467
rect 22385 14433 22419 14467
rect 23673 14433 23707 14467
rect 23857 14433 23891 14467
rect 25329 14433 25363 14467
rect 25513 14433 25547 14467
rect 25973 14433 26007 14467
rect 30757 14433 30791 14467
rect 30941 14433 30975 14467
rect 32229 14433 32263 14467
rect 32413 14433 32447 14467
rect 12541 14365 12575 14399
rect 13185 14365 13219 14399
rect 15485 14365 15519 14399
rect 18153 14365 18187 14399
rect 18337 14365 18371 14399
rect 18889 14365 18923 14399
rect 26249 14365 26283 14399
rect 26709 14365 26743 14399
rect 3341 14297 3375 14331
rect 5365 14297 5399 14331
rect 11529 14297 11563 14331
rect 23213 14297 23247 14331
rect 26065 14297 26099 14331
rect 4445 14229 4479 14263
rect 11989 14229 12023 14263
rect 13553 14229 13587 14263
rect 15025 14229 15059 14263
rect 18245 14229 18279 14263
rect 23765 14229 23799 14263
rect 32321 14229 32355 14263
rect 15301 14025 15335 14059
rect 16221 14025 16255 14059
rect 20821 14025 20855 14059
rect 26617 14025 26651 14059
rect 8309 13957 8343 13991
rect 19349 13957 19383 13991
rect 21557 13957 21591 13991
rect 9229 13889 9263 13923
rect 9413 13889 9447 13923
rect 17969 13889 18003 13923
rect 21005 13889 21039 13923
rect 24409 13889 24443 13923
rect 5457 13821 5491 13855
rect 5825 13821 5859 13855
rect 7021 13821 7055 13855
rect 8125 13821 8159 13855
rect 8309 13821 8343 13855
rect 12265 13821 12299 13855
rect 13001 13821 13035 13855
rect 13921 13821 13955 13855
rect 14105 13821 14139 13855
rect 15485 13821 15519 13855
rect 15577 13821 15611 13855
rect 15705 13821 15739 13855
rect 16221 13821 16255 13855
rect 16405 13821 16439 13855
rect 18236 13821 18270 13855
rect 20729 13821 20763 13855
rect 21465 13821 21499 13855
rect 21649 13821 21683 13855
rect 22661 13821 22695 13855
rect 26525 13821 26559 13855
rect 26709 13821 26743 13855
rect 31217 13821 31251 13855
rect 31953 13821 31987 13855
rect 33057 13821 33091 13855
rect 33241 13821 33275 13855
rect 22937 13753 22971 13787
rect 30941 13753 30975 13787
rect 31769 13753 31803 13787
rect 4031 13685 4065 13719
rect 6929 13685 6963 13719
rect 8769 13685 8803 13719
rect 9137 13685 9171 13719
rect 12541 13685 12575 13719
rect 14289 13685 14323 13719
rect 21005 13685 21039 13719
rect 29469 13685 29503 13719
rect 33425 13685 33459 13719
rect 7757 13481 7791 13515
rect 12357 13481 12391 13515
rect 12725 13481 12759 13515
rect 12817 13481 12851 13515
rect 23029 13481 23063 13515
rect 31309 13481 31343 13515
rect 10333 13413 10367 13447
rect 13737 13413 13771 13447
rect 15025 13413 15059 13447
rect 17233 13413 17267 13447
rect 26985 13413 27019 13447
rect 28825 13413 28859 13447
rect 2881 13345 2915 13379
rect 8585 13345 8619 13379
rect 14749 13345 14783 13379
rect 17325 13345 17359 13379
rect 17601 13345 17635 13379
rect 18245 13345 18279 13379
rect 18429 13345 18463 13379
rect 18797 13345 18831 13379
rect 22753 13345 22787 13379
rect 22845 13345 22879 13379
rect 23857 13345 23891 13379
rect 27169 13345 27203 13379
rect 28641 13345 28675 13379
rect 28917 13345 28951 13379
rect 30665 13345 30699 13379
rect 31217 13345 31251 13379
rect 2973 13277 3007 13311
rect 3157 13277 3191 13311
rect 6009 13277 6043 13311
rect 6285 13277 6319 13311
rect 8309 13277 8343 13311
rect 10057 13277 10091 13311
rect 12909 13277 12943 13311
rect 16773 13277 16807 13311
rect 20085 13277 20119 13311
rect 20361 13277 20395 13311
rect 23029 13277 23063 13311
rect 24133 13277 24167 13311
rect 31861 13277 31895 13311
rect 32137 13277 32171 13311
rect 8493 13209 8527 13243
rect 11805 13209 11839 13243
rect 13553 13209 13587 13243
rect 23949 13209 23983 13243
rect 33609 13209 33643 13243
rect 2513 13141 2547 13175
rect 8401 13141 8435 13175
rect 21833 13141 21867 13175
rect 24041 13141 24075 13175
rect 28457 13141 28491 13175
rect 30573 13141 30607 13175
rect 3203 12937 3237 12971
rect 5365 12937 5399 12971
rect 8677 12937 8711 12971
rect 12633 12937 12667 12971
rect 14013 12937 14047 12971
rect 16313 12937 16347 12971
rect 21649 12937 21683 12971
rect 26065 12937 26099 12971
rect 29561 12937 29595 12971
rect 30297 12937 30331 12971
rect 33057 12937 33091 12971
rect 12357 12869 12391 12903
rect 22753 12869 22787 12903
rect 26157 12869 26191 12903
rect 30389 12869 30423 12903
rect 1777 12801 1811 12835
rect 4721 12801 4755 12835
rect 7941 12801 7975 12835
rect 8125 12801 8159 12835
rect 9137 12801 9171 12835
rect 9321 12801 9355 12835
rect 13185 12801 13219 12835
rect 13829 12801 13863 12835
rect 18705 12801 18739 12835
rect 22569 12801 22603 12835
rect 24041 12801 24075 12835
rect 26249 12801 26283 12835
rect 27813 12801 27847 12835
rect 28089 12801 28123 12835
rect 1409 12733 1443 12767
rect 4905 12733 4939 12767
rect 7849 12733 7883 12767
rect 9045 12733 9079 12767
rect 10057 12733 10091 12767
rect 12173 12733 12207 12767
rect 13001 12733 13035 12767
rect 13093 12733 13127 12767
rect 14105 12733 14139 12767
rect 16221 12733 16255 12767
rect 16405 12733 16439 12767
rect 17693 12733 17727 12767
rect 18061 12733 18095 12767
rect 18521 12733 18555 12767
rect 18797 12733 18831 12767
rect 19165 12733 19199 12767
rect 21833 12733 21867 12767
rect 22845 12733 22879 12767
rect 23765 12733 23799 12767
rect 25973 12733 26007 12767
rect 30113 12733 30147 12767
rect 30205 12733 30239 12767
rect 30481 12733 30515 12767
rect 30941 12733 30975 12767
rect 31125 12733 31159 12767
rect 33057 12733 33091 12767
rect 33333 12733 33367 12767
rect 31309 12665 31343 12699
rect 33241 12665 33275 12699
rect 4997 12597 5031 12631
rect 7481 12597 7515 12631
rect 9873 12597 9907 12631
rect 13829 12597 13863 12631
rect 22569 12597 22603 12631
rect 25513 12597 25547 12631
rect 2789 12393 2823 12427
rect 9505 12393 9539 12427
rect 17693 12393 17727 12427
rect 23581 12393 23615 12427
rect 24133 12393 24167 12427
rect 29561 12393 29595 12427
rect 1777 12325 1811 12359
rect 1961 12325 1995 12359
rect 16865 12325 16899 12359
rect 22753 12325 22787 12359
rect 25881 12325 25915 12359
rect 30481 12325 30515 12359
rect 32321 12325 32355 12359
rect 33609 12325 33643 12359
rect 3157 12257 3191 12291
rect 8585 12257 8619 12291
rect 9873 12257 9907 12291
rect 13093 12257 13127 12291
rect 13277 12257 13311 12291
rect 15393 12257 15427 12291
rect 16773 12257 16807 12291
rect 16957 12257 16991 12291
rect 17601 12257 17635 12291
rect 17785 12257 17819 12291
rect 18797 12257 18831 12291
rect 19993 12257 20027 12291
rect 20177 12257 20211 12291
rect 23029 12257 23063 12291
rect 23489 12257 23523 12291
rect 23673 12257 23707 12291
rect 24133 12257 24167 12291
rect 24317 12257 24351 12291
rect 25237 12257 25271 12291
rect 29377 12257 29411 12291
rect 29561 12257 29595 12291
rect 30757 12257 30791 12291
rect 31033 12257 31067 12291
rect 31125 12257 31159 12291
rect 32137 12257 32171 12291
rect 32413 12257 32447 12291
rect 33425 12257 33459 12291
rect 3065 12189 3099 12223
rect 4629 12189 4663 12223
rect 4997 12189 5031 12223
rect 9965 12189 9999 12223
rect 10057 12189 10091 12223
rect 15669 12189 15703 12223
rect 19073 12189 19107 12223
rect 20085 12189 20119 12223
rect 25605 12189 25639 12223
rect 25421 12121 25455 12155
rect 6423 12053 6457 12087
rect 8493 12053 8527 12087
rect 13277 12053 13311 12087
rect 15485 12053 15519 12087
rect 15577 12053 15611 12087
rect 18889 12053 18923 12087
rect 18981 12053 19015 12087
rect 21281 12053 21315 12087
rect 27353 12053 27387 12087
rect 32137 12053 32171 12087
rect 4997 11849 5031 11883
rect 9137 11849 9171 11883
rect 11069 11849 11103 11883
rect 12909 11849 12943 11883
rect 17417 11849 17451 11883
rect 20361 11849 20395 11883
rect 26525 11849 26559 11883
rect 2881 11781 2915 11815
rect 8585 11781 8619 11815
rect 2697 11713 2731 11747
rect 3525 11713 3559 11747
rect 5457 11713 5491 11747
rect 5549 11713 5583 11747
rect 6837 11713 6871 11747
rect 7113 11713 7147 11747
rect 9781 11713 9815 11747
rect 13553 11713 13587 11747
rect 15853 11713 15887 11747
rect 31401 11713 31435 11747
rect 2973 11645 3007 11679
rect 3433 11645 3467 11679
rect 3617 11645 3651 11679
rect 9505 11645 9539 11679
rect 10517 11645 10551 11679
rect 10977 11645 11011 11679
rect 11161 11645 11195 11679
rect 15586 11645 15620 11679
rect 17509 11645 17543 11679
rect 18981 11645 19015 11679
rect 19237 11645 19271 11679
rect 24409 11645 24443 11679
rect 25053 11645 25087 11679
rect 26433 11645 26467 11679
rect 26617 11645 26651 11679
rect 28181 11645 28215 11679
rect 28457 11645 28491 11679
rect 29561 11645 29595 11679
rect 29745 11645 29779 11679
rect 30757 11645 30791 11679
rect 31125 11645 31159 11679
rect 31493 11645 31527 11679
rect 33149 11645 33183 11679
rect 33333 11645 33367 11679
rect 5365 11577 5399 11611
rect 13277 11577 13311 11611
rect 25789 11577 25823 11611
rect 2697 11509 2731 11543
rect 9597 11509 9631 11543
rect 10425 11509 10459 11543
rect 13369 11509 13403 11543
rect 14473 11509 14507 11543
rect 24317 11509 24351 11543
rect 27997 11509 28031 11543
rect 28365 11509 28399 11543
rect 29653 11509 29687 11543
rect 33333 11509 33367 11543
rect 9505 11305 9539 11339
rect 14912 11305 14946 11339
rect 15761 11305 15795 11339
rect 18061 11305 18095 11339
rect 20637 11305 20671 11339
rect 23213 11305 23247 11339
rect 30573 11305 30607 11339
rect 9689 11237 9723 11271
rect 9873 11237 9907 11271
rect 15117 11237 15151 11271
rect 26065 11237 26099 11271
rect 27813 11237 27847 11271
rect 32137 11237 32171 11271
rect 1409 11169 1443 11203
rect 1777 11169 1811 11203
rect 5273 11169 5307 11203
rect 5365 11169 5399 11203
rect 10425 11169 10459 11203
rect 12725 11169 12759 11203
rect 13553 11169 13587 11203
rect 13737 11169 13771 11203
rect 15669 11169 15703 11203
rect 15853 11169 15887 11203
rect 16957 11169 16991 11203
rect 18061 11169 18095 11203
rect 18245 11169 18279 11203
rect 19073 11169 19107 11203
rect 20453 11169 20487 11203
rect 21741 11169 21775 11203
rect 22385 11169 22419 11203
rect 22569 11169 22603 11203
rect 23029 11169 23063 11203
rect 23581 11169 23615 11203
rect 27077 11169 27111 11203
rect 30481 11169 30515 11203
rect 31309 11169 31343 11203
rect 31861 11169 31895 11203
rect 5457 11101 5491 11135
rect 12173 11101 12207 11135
rect 23857 11101 23891 11135
rect 26157 11101 26191 11135
rect 26249 11101 26283 11135
rect 27537 11101 27571 11135
rect 29285 11101 29319 11135
rect 13553 11033 13587 11067
rect 14749 11033 14783 11067
rect 18981 11033 19015 11067
rect 21833 11033 21867 11067
rect 22477 11033 22511 11067
rect 23673 11033 23707 11067
rect 26985 11033 27019 11067
rect 3203 10965 3237 10999
rect 4905 10965 4939 10999
rect 10682 10965 10716 10999
rect 14933 10965 14967 10999
rect 17233 10965 17267 10999
rect 17417 10965 17451 10999
rect 23765 10965 23799 10999
rect 25697 10965 25731 10999
rect 31217 10965 31251 10999
rect 33609 10965 33643 10999
rect 3341 10761 3375 10795
rect 5779 10761 5813 10795
rect 9781 10761 9815 10795
rect 10425 10761 10459 10795
rect 12081 10761 12115 10795
rect 13369 10761 13403 10795
rect 14381 10761 14415 10795
rect 15301 10761 15335 10795
rect 19809 10761 19843 10795
rect 26893 10761 26927 10795
rect 29193 10761 29227 10795
rect 31769 10761 31803 10795
rect 33149 10761 33183 10795
rect 29423 10693 29457 10727
rect 3985 10625 4019 10659
rect 4353 10625 4387 10659
rect 8861 10625 8895 10659
rect 10977 10625 11011 10659
rect 15485 10625 15519 10659
rect 18613 10625 18647 10659
rect 21189 10625 21223 10659
rect 24409 10625 24443 10659
rect 25145 10625 25179 10659
rect 25421 10625 25455 10659
rect 29285 10625 29319 10659
rect 30757 10625 30791 10659
rect 3433 10557 3467 10591
rect 9689 10557 9723 10591
rect 12265 10557 12299 10591
rect 13001 10557 13035 10591
rect 13277 10557 13311 10591
rect 13461 10557 13495 10591
rect 13921 10557 13955 10591
rect 14197 10557 14231 10591
rect 15209 10557 15243 10591
rect 16221 10557 16255 10591
rect 16405 10557 16439 10591
rect 17601 10557 17635 10591
rect 17877 10557 17911 10591
rect 18245 10557 18279 10591
rect 18705 10557 18739 10591
rect 19257 10557 19291 10591
rect 24142 10557 24176 10591
rect 29101 10557 29135 10591
rect 29561 10557 29595 10591
rect 30665 10557 30699 10591
rect 30941 10557 30975 10591
rect 31125 10557 31159 10591
rect 31585 10557 31619 10591
rect 33057 10557 33091 10591
rect 33241 10557 33275 10591
rect 8585 10489 8619 10523
rect 16313 10489 16347 10523
rect 20922 10489 20956 10523
rect 8217 10421 8251 10455
rect 8677 10421 8711 10455
rect 10793 10421 10827 10455
rect 10885 10421 10919 10455
rect 14013 10421 14047 10455
rect 15485 10421 15519 10455
rect 23029 10421 23063 10455
rect 2789 10217 2823 10251
rect 10241 10217 10275 10251
rect 13277 10217 13311 10251
rect 14749 10217 14783 10251
rect 19993 10217 20027 10251
rect 22201 10217 22235 10251
rect 23949 10217 23983 10251
rect 7389 10149 7423 10183
rect 8493 10149 8527 10183
rect 13645 10149 13679 10183
rect 15862 10149 15896 10183
rect 23213 10149 23247 10183
rect 32597 10149 32631 10183
rect 8217 10081 8251 10115
rect 8309 10081 8343 10115
rect 9505 10081 9539 10115
rect 10425 10081 10459 10115
rect 10517 10081 10551 10115
rect 11345 10081 11379 10115
rect 12909 10081 12943 10115
rect 13461 10081 13495 10115
rect 16129 10081 16163 10115
rect 16681 10081 16715 10115
rect 16957 10081 16991 10115
rect 17417 10081 17451 10115
rect 17785 10081 17819 10115
rect 18153 10081 18187 10115
rect 20177 10081 20211 10115
rect 20269 10081 20303 10115
rect 20821 10081 20855 10115
rect 21088 10081 21122 10115
rect 22661 10081 22695 10115
rect 23305 10081 23339 10115
rect 23857 10081 23891 10115
rect 24041 10081 24075 10115
rect 26617 10081 26651 10115
rect 30757 10081 30791 10115
rect 30849 10081 30883 10115
rect 30941 10081 30975 10115
rect 31125 10081 31159 10115
rect 31585 10081 31619 10115
rect 31769 10081 31803 10115
rect 32413 10081 32447 10115
rect 33241 10081 33275 10115
rect 33425 10081 33459 10115
rect 2881 10013 2915 10047
rect 3065 10013 3099 10047
rect 7481 10013 7515 10047
rect 7665 10013 7699 10047
rect 8493 10013 8527 10047
rect 10241 10013 10275 10047
rect 11437 10013 11471 10047
rect 11529 10013 11563 10047
rect 17693 10013 17727 10047
rect 19993 10013 20027 10047
rect 26893 10013 26927 10047
rect 30481 10013 30515 10047
rect 10977 9945 11011 9979
rect 31861 9945 31895 9979
rect 2421 9877 2455 9911
rect 7021 9877 7055 9911
rect 9597 9877 9631 9911
rect 12725 9877 12759 9911
rect 22845 9877 22879 9911
rect 28365 9877 28399 9911
rect 32781 9877 32815 9911
rect 33333 9877 33367 9911
rect 3203 9673 3237 9707
rect 9137 9673 9171 9707
rect 12081 9673 12115 9707
rect 15669 9673 15703 9707
rect 19809 9673 19843 9707
rect 21373 9673 21407 9707
rect 29929 9673 29963 9707
rect 33241 9673 33275 9707
rect 11069 9605 11103 9639
rect 17601 9605 17635 9639
rect 21465 9605 21499 9639
rect 25973 9605 26007 9639
rect 30757 9605 30791 9639
rect 1777 9537 1811 9571
rect 5549 9537 5583 9571
rect 5641 9537 5675 9571
rect 7113 9537 7147 9571
rect 8585 9537 8619 9571
rect 9781 9537 9815 9571
rect 12725 9537 12759 9571
rect 13829 9537 13863 9571
rect 21281 9537 21315 9571
rect 24593 9537 24627 9571
rect 1409 9469 1443 9503
rect 3893 9469 3927 9503
rect 6837 9469 6871 9503
rect 9505 9469 9539 9503
rect 10333 9469 10367 9503
rect 11161 9469 11195 9503
rect 14473 9469 14507 9503
rect 15577 9469 15611 9503
rect 15761 9469 15795 9503
rect 17325 9469 17359 9503
rect 17601 9469 17635 9503
rect 19717 9469 19751 9503
rect 19901 9469 19935 9503
rect 20637 9469 20671 9503
rect 21557 9469 21591 9503
rect 22569 9469 22603 9503
rect 23857 9469 23891 9503
rect 29009 9469 29043 9503
rect 29469 9469 29503 9503
rect 29745 9469 29779 9503
rect 30849 9469 30883 9503
rect 31217 9469 31251 9503
rect 31401 9469 31435 9503
rect 33057 9469 33091 9503
rect 3709 9401 3743 9435
rect 5457 9401 5491 9435
rect 10425 9401 10459 9435
rect 12449 9401 12483 9435
rect 24838 9401 24872 9435
rect 5089 9333 5123 9367
rect 9597 9333 9631 9367
rect 12541 9333 12575 9367
rect 13277 9333 13311 9367
rect 13645 9333 13679 9367
rect 13737 9333 13771 9367
rect 14565 9333 14599 9367
rect 20821 9333 20855 9367
rect 22661 9333 22695 9367
rect 23765 9333 23799 9367
rect 6055 9129 6089 9163
rect 8493 9129 8527 9163
rect 11437 9129 11471 9163
rect 13645 9129 13679 9163
rect 15761 9129 15795 9163
rect 16497 9129 16531 9163
rect 17233 9129 17267 9163
rect 18245 9129 18279 9163
rect 21557 9129 21591 9163
rect 23581 9129 23615 9163
rect 28917 9129 28951 9163
rect 29469 9129 29503 9163
rect 12725 9061 12759 9095
rect 21465 9061 21499 9095
rect 30757 9061 30791 9095
rect 2789 8993 2823 9027
rect 4629 8993 4663 9027
rect 8401 8993 8435 9027
rect 8585 8993 8619 9027
rect 9505 8993 9539 9027
rect 9689 8993 9723 9027
rect 10517 8993 10551 9027
rect 10701 8993 10735 9027
rect 11345 8993 11379 9027
rect 11529 8993 11563 9027
rect 12633 8993 12667 9027
rect 12817 8993 12851 9027
rect 13277 8993 13311 9027
rect 13461 8993 13495 9027
rect 15853 8993 15887 9027
rect 16313 8993 16347 9027
rect 16497 8993 16531 9027
rect 17141 8993 17175 9027
rect 17325 8993 17359 9027
rect 17785 8993 17819 9027
rect 18797 8993 18831 9027
rect 20729 8993 20763 9027
rect 22661 8993 22695 9027
rect 23857 8993 23891 9027
rect 28733 8993 28767 9027
rect 29377 8993 29411 9027
rect 30941 8993 30975 9027
rect 31125 8993 31159 9027
rect 2697 8925 2731 8959
rect 4261 8925 4295 8959
rect 19073 8925 19107 8959
rect 23581 8925 23615 8959
rect 25697 8925 25731 8959
rect 25973 8925 26007 8959
rect 28457 8925 28491 8959
rect 31585 8925 31619 8959
rect 31861 8925 31895 8959
rect 33609 8925 33643 8959
rect 9597 8857 9631 8891
rect 20545 8857 20579 8891
rect 22845 8857 22879 8891
rect 23765 8857 23799 8891
rect 3065 8789 3099 8823
rect 10701 8789 10735 8823
rect 18061 8789 18095 8823
rect 18889 8789 18923 8823
rect 18981 8789 19015 8823
rect 27445 8789 27479 8823
rect 28549 8789 28583 8823
rect 1593 8585 1627 8619
rect 4445 8585 4479 8619
rect 15945 8585 15979 8619
rect 16313 8585 16347 8619
rect 17325 8585 17359 8619
rect 20085 8585 20119 8619
rect 29745 8585 29779 8619
rect 33057 8585 33091 8619
rect 9413 8517 9447 8551
rect 11253 8517 11287 8551
rect 29101 8517 29135 8551
rect 3341 8449 3375 8483
rect 8861 8449 8895 8483
rect 10609 8449 10643 8483
rect 13185 8449 13219 8483
rect 21281 8449 21315 8483
rect 1409 8381 1443 8415
rect 3157 8381 3191 8415
rect 4261 8381 4295 8415
rect 9597 8381 9631 8415
rect 11437 8381 11471 8415
rect 15209 8381 15243 8415
rect 15393 8381 15427 8415
rect 15853 8381 15887 8415
rect 17509 8381 17543 8415
rect 17969 8381 18003 8415
rect 18705 8381 18739 8415
rect 18972 8381 19006 8415
rect 20821 8381 20855 8415
rect 21465 8381 21499 8415
rect 23305 8381 23339 8415
rect 25145 8381 25179 8415
rect 28181 8381 28215 8415
rect 29285 8381 29319 8415
rect 29975 8381 30009 8415
rect 30113 8381 30147 8415
rect 30205 8381 30239 8415
rect 30389 8381 30423 8415
rect 31401 8381 31435 8415
rect 31585 8381 31619 8415
rect 32045 8381 32079 8415
rect 33333 8381 33367 8415
rect 8585 8313 8619 8347
rect 17877 8313 17911 8347
rect 22569 8313 22603 8347
rect 22753 8313 22787 8347
rect 24878 8313 24912 8347
rect 28273 8313 28307 8347
rect 31493 8313 31527 8347
rect 33057 8313 33091 8347
rect 33241 8313 33275 8347
rect 2789 8245 2823 8279
rect 3249 8245 3283 8279
rect 8217 8245 8251 8279
rect 8677 8245 8711 8279
rect 10057 8245 10091 8279
rect 10425 8245 10459 8279
rect 10517 8245 10551 8279
rect 12633 8245 12667 8279
rect 13001 8245 13035 8279
rect 13093 8245 13127 8279
rect 15393 8245 15427 8279
rect 20637 8245 20671 8279
rect 23489 8245 23523 8279
rect 23765 8245 23799 8279
rect 3203 8041 3237 8075
rect 6331 8041 6365 8075
rect 7757 8041 7791 8075
rect 8125 8041 8159 8075
rect 10425 8041 10459 8075
rect 10885 8041 10919 8075
rect 13093 8041 13127 8075
rect 13461 8041 13495 8075
rect 16129 8041 16163 8075
rect 17693 8041 17727 8075
rect 18245 8041 18279 8075
rect 24133 8041 24167 8075
rect 28733 8041 28767 8075
rect 30481 8041 30515 8075
rect 33517 8041 33551 8075
rect 10793 7973 10827 8007
rect 23305 7973 23339 8007
rect 28089 7973 28123 8007
rect 29561 7973 29595 8007
rect 1409 7905 1443 7939
rect 4537 7905 4571 7939
rect 7021 7905 7055 7939
rect 7113 7905 7147 7939
rect 8217 7905 8251 7939
rect 9965 7905 9999 7939
rect 12081 7905 12115 7939
rect 12173 7905 12207 7939
rect 15016 7905 15050 7939
rect 16773 7905 16807 7939
rect 17417 7905 17451 7939
rect 18337 7905 18371 7939
rect 20545 7905 20579 7939
rect 21640 7905 21674 7939
rect 23397 7905 23431 7939
rect 23857 7905 23891 7939
rect 27813 7905 27847 7939
rect 27997 7905 28031 7939
rect 28641 7905 28675 7939
rect 28825 7905 28859 7939
rect 29285 7905 29319 7939
rect 29377 7905 29411 7939
rect 30757 7905 30791 7939
rect 31309 7905 31343 7939
rect 32321 7905 32355 7939
rect 32873 7905 32907 7939
rect 33333 7905 33367 7939
rect 33609 7905 33643 7939
rect 1777 7837 1811 7871
rect 4905 7837 4939 7871
rect 7300 7837 7334 7871
rect 8401 7837 8435 7871
rect 9689 7837 9723 7871
rect 9873 7837 9907 7871
rect 10977 7837 11011 7871
rect 11897 7837 11931 7871
rect 13553 7837 13587 7871
rect 13645 7837 13679 7871
rect 14749 7837 14783 7871
rect 17693 7837 17727 7871
rect 21373 7837 21407 7871
rect 24133 7837 24167 7871
rect 30665 7837 30699 7871
rect 32413 7837 32447 7871
rect 23949 7769 23983 7803
rect 29561 7769 29595 7803
rect 7205 7701 7239 7735
rect 9781 7701 9815 7735
rect 11989 7701 12023 7735
rect 16681 7701 16715 7735
rect 17509 7701 17543 7735
rect 20453 7701 20487 7735
rect 22753 7701 22787 7735
rect 33333 7701 33367 7735
rect 5181 7497 5215 7531
rect 8493 7497 8527 7531
rect 9045 7497 9079 7531
rect 15669 7497 15703 7531
rect 19717 7497 19751 7531
rect 21465 7497 21499 7531
rect 21557 7497 21591 7531
rect 23305 7497 23339 7531
rect 24133 7497 24167 7531
rect 28917 7497 28951 7531
rect 29929 7497 29963 7531
rect 33241 7497 33275 7531
rect 11069 7429 11103 7463
rect 29009 7429 29043 7463
rect 33425 7429 33459 7463
rect 3157 7361 3191 7395
rect 5641 7361 5675 7395
rect 5733 7361 5767 7395
rect 7849 7361 7883 7395
rect 10241 7361 10275 7395
rect 10425 7361 10459 7395
rect 12633 7361 12667 7395
rect 15577 7361 15611 7395
rect 21649 7361 21683 7395
rect 22661 7361 22695 7395
rect 28917 7361 28951 7395
rect 30665 7361 30699 7395
rect 3065 7293 3099 7327
rect 7573 7293 7607 7327
rect 8585 7293 8619 7327
rect 9045 7293 9079 7327
rect 9229 7293 9263 7327
rect 10149 7293 10183 7327
rect 10977 7293 11011 7327
rect 12449 7293 12483 7327
rect 13645 7293 13679 7327
rect 13829 7293 13863 7327
rect 14473 7293 14507 7327
rect 15761 7293 15795 7327
rect 15853 7293 15887 7327
rect 17325 7293 17359 7327
rect 17581 7293 17615 7327
rect 19625 7293 19659 7327
rect 19809 7293 19843 7327
rect 21373 7293 21407 7327
rect 22569 7293 22603 7327
rect 22753 7293 22787 7327
rect 23213 7293 23247 7327
rect 23397 7293 23431 7327
rect 24041 7293 24075 7327
rect 24225 7293 24259 7327
rect 24685 7293 24719 7327
rect 27997 7293 28031 7327
rect 28181 7293 28215 7327
rect 28273 7293 28307 7327
rect 29101 7293 29135 7327
rect 29837 7293 29871 7327
rect 30021 7293 30055 7327
rect 30573 7293 30607 7327
rect 31217 7293 31251 7327
rect 31309 7293 31343 7327
rect 7665 7225 7699 7259
rect 12541 7225 12575 7259
rect 14565 7225 14599 7259
rect 28733 7225 28767 7259
rect 33057 7225 33091 7259
rect 33273 7225 33307 7259
rect 2605 7157 2639 7191
rect 2973 7157 3007 7191
rect 5549 7157 5583 7191
rect 7205 7157 7239 7191
rect 9781 7157 9815 7191
rect 12081 7157 12115 7191
rect 14013 7157 14047 7191
rect 18705 7157 18739 7191
rect 24869 7157 24903 7191
rect 27813 7157 27847 7191
rect 10701 6953 10735 6987
rect 12817 6953 12851 6987
rect 17877 6953 17911 6987
rect 27905 6953 27939 6987
rect 33609 6953 33643 6987
rect 5273 6885 5307 6919
rect 11069 6885 11103 6919
rect 13737 6885 13771 6919
rect 1869 6817 1903 6851
rect 5365 6817 5399 6851
rect 11989 6817 12023 6851
rect 12725 6817 12759 6851
rect 12909 6817 12943 6851
rect 13369 6817 13403 6851
rect 13553 6817 13587 6851
rect 15761 6817 15795 6851
rect 16681 6817 16715 6851
rect 16773 6817 16807 6851
rect 17877 6817 17911 6851
rect 18061 6817 18095 6851
rect 19073 6817 19107 6851
rect 20637 6817 20671 6851
rect 21189 6817 21223 6851
rect 21281 6817 21315 6851
rect 21925 6817 21959 6851
rect 23765 6817 23799 6851
rect 25605 6817 25639 6851
rect 27813 6817 27847 6851
rect 28733 6817 28767 6851
rect 28917 6817 28951 6851
rect 29377 6817 29411 6851
rect 29561 6817 29595 6851
rect 1501 6749 1535 6783
rect 5457 6749 5491 6783
rect 11161 6749 11195 6783
rect 11253 6749 11287 6783
rect 15485 6749 15519 6783
rect 18797 6749 18831 6783
rect 20361 6749 20395 6783
rect 23857 6749 23891 6783
rect 24041 6749 24075 6783
rect 25881 6749 25915 6783
rect 27353 6749 27387 6783
rect 29469 6749 29503 6783
rect 31861 6749 31895 6783
rect 32137 6749 32171 6783
rect 20545 6681 20579 6715
rect 3295 6613 3329 6647
rect 4905 6613 4939 6647
rect 12173 6613 12207 6647
rect 15577 6613 15611 6647
rect 15669 6613 15703 6647
rect 18889 6613 18923 6647
rect 18981 6613 19015 6647
rect 20453 6613 20487 6647
rect 21741 6613 21775 6647
rect 23949 6613 23983 6647
rect 28825 6613 28859 6647
rect 5687 6409 5721 6443
rect 9413 6409 9447 6443
rect 10977 6409 11011 6443
rect 13369 6409 13403 6443
rect 16221 6409 16255 6443
rect 22753 6409 22787 6443
rect 29285 6409 29319 6443
rect 30021 6409 30055 6443
rect 30205 6409 30239 6443
rect 33241 6409 33275 6443
rect 12817 6341 12851 6375
rect 4261 6273 4295 6307
rect 6929 6273 6963 6307
rect 7205 6273 7239 6307
rect 10057 6273 10091 6307
rect 13829 6273 13863 6307
rect 13921 6273 13955 6307
rect 14841 6273 14875 6307
rect 19533 6273 19567 6307
rect 19993 6273 20027 6307
rect 22569 6273 22603 6307
rect 29193 6273 29227 6307
rect 3893 6205 3927 6239
rect 10885 6205 10919 6239
rect 12725 6205 12759 6239
rect 12909 6205 12943 6239
rect 13737 6205 13771 6239
rect 15108 6205 15142 6239
rect 19266 6205 19300 6239
rect 20260 6205 20294 6239
rect 22845 6205 22879 6239
rect 23765 6205 23799 6239
rect 23857 6205 23891 6239
rect 24317 6205 24351 6239
rect 24573 6205 24607 6239
rect 28089 6205 28123 6239
rect 28273 6205 28307 6239
rect 28365 6205 28399 6239
rect 29377 6205 29411 6239
rect 29469 6205 29503 6239
rect 30849 6205 30883 6239
rect 31493 6205 31527 6239
rect 33057 6205 33091 6239
rect 33241 6205 33275 6239
rect 8953 6137 8987 6171
rect 9873 6137 9907 6171
rect 30173 6137 30207 6171
rect 30389 6137 30423 6171
rect 9781 6069 9815 6103
rect 18153 6069 18187 6103
rect 21373 6069 21407 6103
rect 22569 6069 22603 6103
rect 25697 6069 25731 6103
rect 27905 6069 27939 6103
rect 30941 6069 30975 6103
rect 31585 6069 31619 6103
rect 2973 5865 3007 5899
rect 5687 5865 5721 5899
rect 8217 5865 8251 5899
rect 10517 5865 10551 5899
rect 15945 5865 15979 5899
rect 16497 5865 16531 5899
rect 20085 5865 20119 5899
rect 20637 5865 20671 5899
rect 29285 5865 29319 5899
rect 8401 5797 8435 5831
rect 11805 5797 11839 5831
rect 22376 5797 22410 5831
rect 27813 5797 27847 5831
rect 30941 5797 30975 5831
rect 8585 5729 8619 5763
rect 9781 5729 9815 5763
rect 10149 5729 10183 5763
rect 10425 5729 10459 5763
rect 16037 5729 16071 5763
rect 16497 5729 16531 5763
rect 16681 5729 16715 5763
rect 17325 5729 17359 5763
rect 17417 5729 17451 5763
rect 18245 5729 18279 5763
rect 19993 5729 20027 5763
rect 20177 5729 20211 5763
rect 20637 5729 20671 5763
rect 20821 5729 20855 5763
rect 24133 5729 24167 5763
rect 3065 5661 3099 5695
rect 3249 5661 3283 5695
rect 7113 5661 7147 5695
rect 7481 5661 7515 5695
rect 11529 5661 11563 5695
rect 17601 5661 17635 5695
rect 22109 5661 22143 5695
rect 25329 5661 25363 5695
rect 25605 5661 25639 5695
rect 27537 5661 27571 5695
rect 31861 5661 31895 5695
rect 32137 5661 32171 5695
rect 17509 5593 17543 5627
rect 24041 5593 24075 5627
rect 2605 5525 2639 5559
rect 13277 5525 13311 5559
rect 18153 5525 18187 5559
rect 23489 5525 23523 5559
rect 27077 5525 27111 5559
rect 31033 5525 31067 5559
rect 33609 5525 33643 5559
rect 3203 5321 3237 5355
rect 5917 5321 5951 5355
rect 9137 5321 9171 5355
rect 10609 5321 10643 5355
rect 13461 5321 13495 5355
rect 20729 5321 20763 5355
rect 22661 5321 22695 5355
rect 23305 5321 23339 5355
rect 24225 5321 24259 5355
rect 25513 5321 25547 5355
rect 31953 5321 31987 5355
rect 30941 5253 30975 5287
rect 1409 5185 1443 5219
rect 1777 5185 1811 5219
rect 5365 5185 5399 5219
rect 5457 5185 5491 5219
rect 9505 5185 9539 5219
rect 10333 5185 10367 5219
rect 16129 5185 16163 5219
rect 17325 5185 17359 5219
rect 20913 5185 20947 5219
rect 25973 5185 26007 5219
rect 26065 5185 26099 5219
rect 9321 5117 9355 5151
rect 9597 5117 9631 5151
rect 10241 5117 10275 5151
rect 13369 5117 13403 5151
rect 17581 5117 17615 5151
rect 20637 5117 20671 5151
rect 21373 5117 21407 5151
rect 22753 5117 22787 5151
rect 23213 5117 23247 5151
rect 23397 5117 23431 5151
rect 24133 5117 24167 5151
rect 24317 5117 24351 5151
rect 30205 5117 30239 5151
rect 30389 5117 30423 5151
rect 31033 5117 31067 5151
rect 31217 5117 31251 5151
rect 31677 5117 31711 5151
rect 31953 5117 31987 5151
rect 33425 5117 33459 5151
rect 15853 5049 15887 5083
rect 21465 5049 21499 5083
rect 5549 4981 5583 5015
rect 15485 4981 15519 5015
rect 15945 4981 15979 5015
rect 18705 4981 18739 5015
rect 20913 4981 20947 5015
rect 25881 4981 25915 5015
rect 30297 4981 30331 5015
rect 31769 4981 31803 5015
rect 33517 4981 33551 5015
rect 17785 4777 17819 4811
rect 22385 4777 22419 4811
rect 23305 4777 23339 4811
rect 31953 4777 31987 4811
rect 1961 4709 1995 4743
rect 2973 4709 3007 4743
rect 15025 4709 15059 4743
rect 21250 4709 21284 4743
rect 30665 4709 30699 4743
rect 31309 4709 31343 4743
rect 33425 4709 33459 4743
rect 33609 4709 33643 4743
rect 4261 4641 4295 4675
rect 14749 4641 14783 4675
rect 17785 4641 17819 4675
rect 17969 4641 18003 4675
rect 18797 4641 18831 4675
rect 18889 4641 18923 4675
rect 19993 4641 20027 4675
rect 20177 4641 20211 4675
rect 23213 4641 23247 4675
rect 27445 4641 27479 4675
rect 27629 4641 27663 4675
rect 27721 4641 27755 4675
rect 30573 4641 30607 4675
rect 30757 4641 30791 4675
rect 31217 4641 31251 4675
rect 31493 4641 31527 4675
rect 31953 4641 31987 4675
rect 32137 4641 32171 4675
rect 3065 4573 3099 4607
rect 3249 4573 3283 4607
rect 4629 4573 4663 4607
rect 19073 4573 19107 4607
rect 20085 4573 20119 4607
rect 21005 4573 21039 4607
rect 23397 4573 23431 4607
rect 1869 4437 1903 4471
rect 2605 4437 2639 4471
rect 6055 4437 6089 4471
rect 16497 4437 16531 4471
rect 18981 4437 19015 4471
rect 22845 4437 22879 4471
rect 27261 4437 27295 4471
rect 31493 4437 31527 4471
rect 3755 4233 3789 4267
rect 9584 4233 9618 4267
rect 14491 4233 14525 4267
rect 20913 4233 20947 4267
rect 22924 4233 22958 4267
rect 28089 4233 28123 4267
rect 31401 4233 31435 4267
rect 1961 4097 1995 4131
rect 2329 4097 2363 4131
rect 5365 4097 5399 4131
rect 5457 4097 5491 4131
rect 9321 4097 9355 4131
rect 11069 4097 11103 4131
rect 13001 4097 13035 4131
rect 14749 4097 14783 4131
rect 18889 4097 18923 4131
rect 28457 4097 28491 4131
rect 30665 4097 30699 4131
rect 31493 4097 31527 4131
rect 19145 4029 19179 4063
rect 20821 4029 20855 4063
rect 21005 4029 21039 4063
rect 22661 4029 22695 4063
rect 28365 4029 28399 4063
rect 29193 4029 29227 4063
rect 29469 4029 29503 4063
rect 30297 4029 30331 4063
rect 30481 4029 30515 4063
rect 31217 4029 31251 4063
rect 31309 4029 31343 4063
rect 5549 3961 5583 3995
rect 5917 3893 5951 3927
rect 20269 3893 20303 3927
rect 24409 3893 24443 3927
rect 29009 3893 29043 3927
rect 29377 3893 29411 3927
rect 4261 3689 4295 3723
rect 5595 3689 5629 3723
rect 29561 3689 29595 3723
rect 33333 3689 33367 3723
rect 26801 3621 26835 3655
rect 28549 3621 28583 3655
rect 31861 3621 31895 3655
rect 4629 3553 4663 3587
rect 4721 3553 4755 3587
rect 7021 3553 7055 3587
rect 7389 3553 7423 3587
rect 17253 3553 17287 3587
rect 17509 3553 17543 3587
rect 18153 3553 18187 3587
rect 18245 3553 18279 3587
rect 21005 3553 21039 3587
rect 29285 3553 29319 3587
rect 29377 3553 29411 3587
rect 30757 3553 30791 3587
rect 31585 3553 31619 3587
rect 4905 3485 4939 3519
rect 18429 3485 18463 3519
rect 26525 3485 26559 3519
rect 29561 3485 29595 3519
rect 30481 3485 30515 3519
rect 30573 3417 30607 3451
rect 16129 3349 16163 3383
rect 18337 3349 18371 3383
rect 20913 3349 20947 3383
rect 30665 3349 30699 3383
rect 17509 3145 17543 3179
rect 20545 3145 20579 3179
rect 30205 3145 30239 3179
rect 30757 3145 30791 3179
rect 17417 3009 17451 3043
rect 17601 3009 17635 3043
rect 20729 3009 20763 3043
rect 21281 3009 21315 3043
rect 28457 3009 28491 3043
rect 28733 3009 28767 3043
rect 17325 2941 17359 2975
rect 18061 2941 18095 2975
rect 18328 2941 18362 2975
rect 20453 2941 20487 2975
rect 21189 2941 21223 2975
rect 21373 2941 21407 2975
rect 30665 2941 30699 2975
rect 19441 2805 19475 2839
rect 20729 2805 20763 2839
rect 5733 2601 5767 2635
rect 13829 2601 13863 2635
rect 17693 2601 17727 2635
rect 18429 2601 18463 2635
rect 21925 2601 21959 2635
rect 1961 2533 1995 2567
rect 11253 2533 11287 2567
rect 16497 2533 16531 2567
rect 19165 2533 19199 2567
rect 20790 2533 20824 2567
rect 23121 2533 23155 2567
rect 25789 2533 25823 2567
rect 28457 2533 28491 2567
rect 31125 2533 31159 2567
rect 31769 2533 31803 2567
rect 32505 2533 32539 2567
rect 2881 2465 2915 2499
rect 5549 2465 5583 2499
rect 8493 2465 8527 2499
rect 14013 2465 14047 2499
rect 17601 2465 17635 2499
rect 17785 2465 17819 2499
rect 18429 2465 18463 2499
rect 18613 2465 18647 2499
rect 20545 2465 20579 2499
rect 3065 2397 3099 2431
rect 1777 2329 1811 2363
rect 8309 2329 8343 2363
rect 11069 2329 11103 2363
rect 19349 2329 19383 2363
rect 22937 2329 22971 2363
rect 25605 2329 25639 2363
rect 28273 2329 28307 2363
rect 30941 2329 30975 2363
rect 31953 2329 31987 2363
rect 32689 2329 32723 2363
rect 16589 2261 16623 2295
<< metal1 >>
rect 7098 35436 7104 35488
rect 7156 35476 7162 35488
rect 15838 35476 15844 35488
rect 7156 35448 15844 35476
rect 7156 35436 7162 35448
rect 15838 35436 15844 35448
rect 15896 35436 15902 35488
rect 1104 35386 34316 35408
rect 1104 35334 12052 35386
rect 12104 35334 12116 35386
rect 12168 35334 12180 35386
rect 12232 35334 12244 35386
rect 12296 35334 23123 35386
rect 23175 35334 23187 35386
rect 23239 35334 23251 35386
rect 23303 35334 23315 35386
rect 23367 35334 34316 35386
rect 1104 35312 34316 35334
rect 1581 35275 1639 35281
rect 1581 35241 1593 35275
rect 1627 35272 1639 35275
rect 7098 35272 7104 35284
rect 1627 35244 7104 35272
rect 1627 35241 1639 35244
rect 1581 35235 1639 35241
rect 7098 35232 7104 35244
rect 7156 35232 7162 35284
rect 7193 35275 7251 35281
rect 7193 35241 7205 35275
rect 7239 35272 7251 35275
rect 12618 35272 12624 35284
rect 7239 35244 12624 35272
rect 7239 35241 7251 35244
rect 7193 35235 7251 35241
rect 12618 35232 12624 35244
rect 12676 35232 12682 35284
rect 21634 35232 21640 35284
rect 21692 35272 21698 35284
rect 21729 35275 21787 35281
rect 21729 35272 21741 35275
rect 21692 35244 21741 35272
rect 21692 35232 21698 35244
rect 21729 35241 21741 35244
rect 21775 35241 21787 35275
rect 21729 35235 21787 35241
rect 24394 35232 24400 35284
rect 24452 35272 24458 35284
rect 24489 35275 24547 35281
rect 24489 35272 24501 35275
rect 24452 35244 24501 35272
rect 24452 35232 24458 35244
rect 24489 35241 24501 35244
rect 24535 35241 24547 35275
rect 24489 35235 24547 35241
rect 10594 35204 10600 35216
rect 8036 35176 10456 35204
rect 10555 35176 10600 35204
rect 1394 35136 1400 35148
rect 1355 35108 1400 35136
rect 1394 35096 1400 35108
rect 1452 35096 1458 35148
rect 2774 35136 2780 35148
rect 2735 35108 2780 35136
rect 2774 35096 2780 35108
rect 2832 35096 2838 35148
rect 5074 35136 5080 35148
rect 5035 35108 5080 35136
rect 5074 35096 5080 35108
rect 5132 35096 5138 35148
rect 7377 35139 7435 35145
rect 7377 35105 7389 35139
rect 7423 35136 7435 35139
rect 7834 35136 7840 35148
rect 7423 35108 7840 35136
rect 7423 35105 7435 35108
rect 7377 35099 7435 35105
rect 7834 35096 7840 35108
rect 7892 35096 7898 35148
rect 8036 35077 8064 35176
rect 8205 35139 8263 35145
rect 8205 35105 8217 35139
rect 8251 35136 8263 35139
rect 8386 35136 8392 35148
rect 8251 35108 8392 35136
rect 8251 35105 8263 35108
rect 8205 35099 8263 35105
rect 8386 35096 8392 35108
rect 8444 35096 8450 35148
rect 8021 35071 8079 35077
rect 8021 35037 8033 35071
rect 8067 35037 8079 35071
rect 8021 35031 8079 35037
rect 8113 35071 8171 35077
rect 8113 35037 8125 35071
rect 8159 35037 8171 35071
rect 8113 35031 8171 35037
rect 5261 35003 5319 35009
rect 5261 34969 5273 35003
rect 5307 35000 5319 35003
rect 8128 35000 8156 35031
rect 8202 35000 8208 35012
rect 5307 34972 8064 35000
rect 8128 34972 8208 35000
rect 5307 34969 5319 34972
rect 5261 34963 5319 34969
rect 2958 34932 2964 34944
rect 2919 34904 2964 34932
rect 2958 34892 2964 34904
rect 3016 34892 3022 34944
rect 8036 34932 8064 34972
rect 8202 34960 8208 34972
rect 8260 34960 8266 35012
rect 10428 35000 10456 35176
rect 10594 35164 10600 35176
rect 10652 35164 10658 35216
rect 13354 35204 13360 35216
rect 13315 35176 13360 35204
rect 13354 35164 13360 35176
rect 13412 35164 13418 35216
rect 13446 35164 13452 35216
rect 13504 35204 13510 35216
rect 27062 35204 27068 35216
rect 13504 35176 27068 35204
rect 13504 35164 13510 35176
rect 27062 35164 27068 35176
rect 27120 35164 27126 35216
rect 27154 35164 27160 35216
rect 27212 35164 27218 35216
rect 32585 35207 32643 35213
rect 32585 35173 32597 35207
rect 32631 35204 32643 35207
rect 32674 35204 32680 35216
rect 32631 35176 32680 35204
rect 32631 35173 32643 35176
rect 32585 35167 32643 35173
rect 32674 35164 32680 35176
rect 32732 35164 32738 35216
rect 10781 35139 10839 35145
rect 10781 35105 10793 35139
rect 10827 35105 10839 35139
rect 10781 35099 10839 35105
rect 13541 35139 13599 35145
rect 13541 35105 13553 35139
rect 13587 35136 13599 35139
rect 14458 35136 14464 35148
rect 13587 35108 14464 35136
rect 13587 35105 13599 35108
rect 13541 35099 13599 35105
rect 10796 35068 10824 35099
rect 14458 35096 14464 35108
rect 14516 35096 14522 35148
rect 16114 35096 16120 35148
rect 16172 35136 16178 35148
rect 16301 35139 16359 35145
rect 16301 35136 16313 35139
rect 16172 35108 16313 35136
rect 16172 35096 16178 35108
rect 16301 35105 16313 35108
rect 16347 35105 16359 35139
rect 18874 35136 18880 35148
rect 18835 35108 18880 35136
rect 16301 35099 16359 35105
rect 18874 35096 18880 35108
rect 18932 35096 18938 35148
rect 21818 35136 21824 35148
rect 21779 35108 21824 35136
rect 21818 35096 21824 35108
rect 21876 35096 21882 35148
rect 24581 35139 24639 35145
rect 24581 35105 24593 35139
rect 24627 35105 24639 35139
rect 27172 35136 27200 35164
rect 27341 35139 27399 35145
rect 27341 35136 27353 35139
rect 27172 35108 27353 35136
rect 24581 35099 24639 35105
rect 27341 35105 27353 35108
rect 27387 35105 27399 35139
rect 27341 35099 27399 35105
rect 14274 35068 14280 35080
rect 10796 35040 14280 35068
rect 14274 35028 14280 35040
rect 14332 35028 14338 35080
rect 20070 35028 20076 35080
rect 20128 35068 20134 35080
rect 24596 35068 24624 35099
rect 29914 35096 29920 35148
rect 29972 35136 29978 35148
rect 30009 35139 30067 35145
rect 30009 35136 30021 35139
rect 29972 35108 30021 35136
rect 29972 35096 29978 35108
rect 30009 35105 30021 35108
rect 30055 35105 30067 35139
rect 30009 35099 30067 35105
rect 31941 35139 31999 35145
rect 31941 35105 31953 35139
rect 31987 35136 31999 35139
rect 34974 35136 34980 35148
rect 31987 35108 34980 35136
rect 31987 35105 31999 35108
rect 31941 35099 31999 35105
rect 34974 35096 34980 35108
rect 35032 35096 35038 35148
rect 20128 35040 24624 35068
rect 27157 35071 27215 35077
rect 20128 35028 20134 35040
rect 27157 35037 27169 35071
rect 27203 35068 27215 35071
rect 29270 35068 29276 35080
rect 27203 35040 29276 35068
rect 27203 35037 27215 35040
rect 27157 35031 27215 35037
rect 29270 35028 29276 35040
rect 29328 35028 29334 35080
rect 12526 35000 12532 35012
rect 10428 34972 12532 35000
rect 12526 34960 12532 34972
rect 12584 34960 12590 35012
rect 8478 34932 8484 34944
rect 8036 34904 8484 34932
rect 8478 34892 8484 34904
rect 8536 34892 8542 34944
rect 8573 34935 8631 34941
rect 8573 34901 8585 34935
rect 8619 34932 8631 34935
rect 8662 34932 8668 34944
rect 8619 34904 8668 34932
rect 8619 34901 8631 34904
rect 8573 34895 8631 34901
rect 8662 34892 8668 34904
rect 8720 34892 8726 34944
rect 15286 34892 15292 34944
rect 15344 34932 15350 34944
rect 16117 34935 16175 34941
rect 16117 34932 16129 34935
rect 15344 34904 16129 34932
rect 15344 34892 15350 34904
rect 16117 34901 16129 34904
rect 16163 34901 16175 34935
rect 16117 34895 16175 34901
rect 18874 34892 18880 34944
rect 18932 34932 18938 34944
rect 19061 34935 19119 34941
rect 19061 34932 19073 34935
rect 18932 34904 19073 34932
rect 18932 34892 18938 34904
rect 19061 34901 19073 34904
rect 19107 34901 19119 34935
rect 19061 34895 19119 34901
rect 29454 34892 29460 34944
rect 29512 34932 29518 34944
rect 29825 34935 29883 34941
rect 29825 34932 29837 34935
rect 29512 34904 29837 34932
rect 29512 34892 29518 34904
rect 29825 34901 29837 34904
rect 29871 34901 29883 34935
rect 29825 34895 29883 34901
rect 31757 34935 31815 34941
rect 31757 34901 31769 34935
rect 31803 34932 31815 34935
rect 32306 34932 32312 34944
rect 31803 34904 32312 34932
rect 31803 34901 31815 34904
rect 31757 34895 31815 34901
rect 32306 34892 32312 34904
rect 32364 34892 32370 34944
rect 32490 34932 32496 34944
rect 32451 34904 32496 34932
rect 32490 34892 32496 34904
rect 32548 34892 32554 34944
rect 1104 34842 34316 34864
rect 1104 34790 6517 34842
rect 6569 34790 6581 34842
rect 6633 34790 6645 34842
rect 6697 34790 6709 34842
rect 6761 34790 17588 34842
rect 17640 34790 17652 34842
rect 17704 34790 17716 34842
rect 17768 34790 17780 34842
rect 17832 34790 28658 34842
rect 28710 34790 28722 34842
rect 28774 34790 28786 34842
rect 28838 34790 28850 34842
rect 28902 34790 34316 34842
rect 1104 34768 34316 34790
rect 8386 34728 8392 34740
rect 8347 34700 8392 34728
rect 8386 34688 8392 34700
rect 8444 34688 8450 34740
rect 8478 34688 8484 34740
rect 8536 34728 8542 34740
rect 8536 34700 12756 34728
rect 8536 34688 8542 34700
rect 2958 34620 2964 34672
rect 3016 34660 3022 34672
rect 3016 34632 7972 34660
rect 3016 34620 3022 34632
rect 7190 34552 7196 34604
rect 7248 34592 7254 34604
rect 7944 34601 7972 34632
rect 9674 34620 9680 34672
rect 9732 34660 9738 34672
rect 9815 34663 9873 34669
rect 9815 34660 9827 34663
rect 9732 34632 9827 34660
rect 9732 34620 9738 34632
rect 9815 34629 9827 34632
rect 9861 34629 9873 34663
rect 9815 34623 9873 34629
rect 12069 34663 12127 34669
rect 12069 34629 12081 34663
rect 12115 34629 12127 34663
rect 12069 34623 12127 34629
rect 7745 34595 7803 34601
rect 7745 34592 7757 34595
rect 7248 34564 7757 34592
rect 7248 34552 7254 34564
rect 7745 34561 7757 34564
rect 7791 34561 7803 34595
rect 7745 34555 7803 34561
rect 7929 34595 7987 34601
rect 7929 34561 7941 34595
rect 7975 34561 7987 34595
rect 12084 34592 12112 34623
rect 7929 34555 7987 34561
rect 9692 34564 12112 34592
rect 9692 34533 9720 34564
rect 12526 34552 12532 34604
rect 12584 34592 12590 34604
rect 12621 34595 12679 34601
rect 12621 34592 12633 34595
rect 12584 34564 12633 34592
rect 12584 34552 12590 34564
rect 12621 34561 12633 34564
rect 12667 34561 12679 34595
rect 12728 34592 12756 34700
rect 27062 34688 27068 34740
rect 27120 34728 27126 34740
rect 29365 34731 29423 34737
rect 29365 34728 29377 34731
rect 27120 34700 29377 34728
rect 27120 34688 27126 34700
rect 29365 34697 29377 34700
rect 29411 34697 29423 34731
rect 29365 34691 29423 34697
rect 15197 34663 15255 34669
rect 15197 34629 15209 34663
rect 15243 34660 15255 34663
rect 16390 34660 16396 34672
rect 15243 34632 16396 34660
rect 15243 34629 15255 34632
rect 15197 34623 15255 34629
rect 16390 34620 16396 34632
rect 16448 34620 16454 34672
rect 12728 34564 13952 34592
rect 12621 34555 12679 34561
rect 9677 34527 9735 34533
rect 9677 34493 9689 34527
rect 9723 34493 9735 34527
rect 9950 34524 9956 34536
rect 9911 34496 9956 34524
rect 9677 34487 9735 34493
rect 9950 34484 9956 34496
rect 10008 34484 10014 34536
rect 10137 34527 10195 34533
rect 10137 34493 10149 34527
rect 10183 34524 10195 34527
rect 10502 34524 10508 34536
rect 10183 34496 10508 34524
rect 10183 34493 10195 34496
rect 10137 34487 10195 34493
rect 10502 34484 10508 34496
rect 10560 34484 10566 34536
rect 12636 34524 12664 34555
rect 12986 34524 12992 34536
rect 12636 34496 12992 34524
rect 12986 34484 12992 34496
rect 13044 34484 13050 34536
rect 13814 34524 13820 34536
rect 13775 34496 13820 34524
rect 13814 34484 13820 34496
rect 13872 34484 13878 34536
rect 13924 34524 13952 34564
rect 19886 34552 19892 34604
rect 19944 34592 19950 34604
rect 20855 34595 20913 34601
rect 20855 34592 20867 34595
rect 19944 34564 20867 34592
rect 19944 34552 19950 34564
rect 20855 34561 20867 34564
rect 20901 34561 20913 34595
rect 20855 34555 20913 34561
rect 14073 34527 14131 34533
rect 14073 34524 14085 34527
rect 13924 34496 14085 34524
rect 14073 34493 14085 34496
rect 14119 34493 14131 34527
rect 14073 34487 14131 34493
rect 17126 34484 17132 34536
rect 17184 34524 17190 34536
rect 19061 34527 19119 34533
rect 19061 34524 19073 34527
rect 17184 34496 19073 34524
rect 17184 34484 17190 34496
rect 19061 34493 19073 34496
rect 19107 34493 19119 34527
rect 19426 34524 19432 34536
rect 19387 34496 19432 34524
rect 19061 34487 19119 34493
rect 19426 34484 19432 34496
rect 19484 34484 19490 34536
rect 22649 34527 22707 34533
rect 22649 34493 22661 34527
rect 22695 34493 22707 34527
rect 23014 34524 23020 34536
rect 22975 34496 23020 34524
rect 22649 34487 22707 34493
rect 8021 34391 8079 34397
rect 8021 34357 8033 34391
rect 8067 34388 8079 34391
rect 8202 34388 8208 34400
rect 8067 34360 8208 34388
rect 8067 34357 8079 34360
rect 8021 34351 8079 34357
rect 8202 34348 8208 34360
rect 8260 34348 8266 34400
rect 10134 34388 10140 34400
rect 10095 34360 10140 34388
rect 10134 34348 10140 34360
rect 10192 34348 10198 34400
rect 12434 34388 12440 34400
rect 12395 34360 12440 34388
rect 12434 34348 12440 34360
rect 12492 34348 12498 34400
rect 12526 34348 12532 34400
rect 12584 34388 12590 34400
rect 20456 34388 20484 34442
rect 20990 34416 20996 34468
rect 21048 34456 21054 34468
rect 22664 34456 22692 34487
rect 23014 34484 23020 34496
rect 23072 34484 23078 34536
rect 29454 34524 29460 34536
rect 29415 34496 29460 34524
rect 29454 34484 29460 34496
rect 29512 34484 29518 34536
rect 21048 34428 22692 34456
rect 21048 34416 21054 34428
rect 20714 34388 20720 34400
rect 12584 34360 12629 34388
rect 20456 34360 20720 34388
rect 12584 34348 12590 34360
rect 20714 34348 20720 34360
rect 20772 34388 20778 34400
rect 21910 34388 21916 34400
rect 20772 34360 21916 34388
rect 20772 34348 20778 34360
rect 21910 34348 21916 34360
rect 21968 34388 21974 34400
rect 23400 34388 23428 34442
rect 21968 34360 23428 34388
rect 21968 34348 21974 34360
rect 23750 34348 23756 34400
rect 23808 34388 23814 34400
rect 24443 34391 24501 34397
rect 24443 34388 24455 34391
rect 23808 34360 24455 34388
rect 23808 34348 23814 34360
rect 24443 34357 24455 34360
rect 24489 34357 24501 34391
rect 24443 34351 24501 34357
rect 1104 34298 34316 34320
rect 1104 34246 12052 34298
rect 12104 34246 12116 34298
rect 12168 34246 12180 34298
rect 12232 34246 12244 34298
rect 12296 34246 23123 34298
rect 23175 34246 23187 34298
rect 23239 34246 23251 34298
rect 23303 34246 23315 34298
rect 23367 34246 34316 34298
rect 1104 34224 34316 34246
rect 12253 34187 12311 34193
rect 12253 34153 12265 34187
rect 12299 34184 12311 34187
rect 12434 34184 12440 34196
rect 12299 34156 12440 34184
rect 12299 34153 12311 34156
rect 12253 34147 12311 34153
rect 12434 34144 12440 34156
rect 12492 34144 12498 34196
rect 12526 34144 12532 34196
rect 12584 34184 12590 34196
rect 12621 34187 12679 34193
rect 12621 34184 12633 34187
rect 12584 34156 12633 34184
rect 12584 34144 12590 34156
rect 12621 34153 12633 34156
rect 12667 34153 12679 34187
rect 12621 34147 12679 34153
rect 12713 34187 12771 34193
rect 12713 34153 12725 34187
rect 12759 34184 12771 34187
rect 13446 34184 13452 34196
rect 12759 34156 13452 34184
rect 12759 34153 12771 34156
rect 12713 34147 12771 34153
rect 13446 34144 13452 34156
rect 13504 34144 13510 34196
rect 23014 34144 23020 34196
rect 23072 34184 23078 34196
rect 23293 34187 23351 34193
rect 23293 34184 23305 34187
rect 23072 34156 23305 34184
rect 23072 34144 23078 34156
rect 23293 34153 23305 34156
rect 23339 34153 23351 34187
rect 23750 34184 23756 34196
rect 23711 34156 23756 34184
rect 23293 34147 23351 34153
rect 23750 34144 23756 34156
rect 23808 34144 23814 34196
rect 10134 34125 10140 34128
rect 10128 34116 10140 34125
rect 10095 34088 10140 34116
rect 10128 34079 10140 34088
rect 10134 34076 10140 34079
rect 10192 34076 10198 34128
rect 20714 34116 20720 34128
rect 18538 34102 20720 34116
rect 18524 34088 20720 34102
rect 13446 34048 13452 34060
rect 13407 34020 13452 34048
rect 13446 34008 13452 34020
rect 13504 34008 13510 34060
rect 13814 34008 13820 34060
rect 13872 34048 13878 34060
rect 16298 34048 16304 34060
rect 13872 34020 16304 34048
rect 13872 34008 13878 34020
rect 16298 34008 16304 34020
rect 16356 34048 16362 34060
rect 17126 34048 17132 34060
rect 16356 34020 17132 34048
rect 16356 34008 16362 34020
rect 17126 34008 17132 34020
rect 17184 34008 17190 34060
rect 9674 33940 9680 33992
rect 9732 33980 9738 33992
rect 9861 33983 9919 33989
rect 9861 33980 9873 33983
rect 9732 33952 9873 33980
rect 9732 33940 9738 33952
rect 9861 33949 9873 33952
rect 9907 33949 9919 33983
rect 12802 33980 12808 33992
rect 12763 33952 12808 33980
rect 9861 33943 9919 33949
rect 12802 33940 12808 33952
rect 12860 33940 12866 33992
rect 17497 33983 17555 33989
rect 17497 33949 17509 33983
rect 17543 33980 17555 33983
rect 18046 33980 18052 33992
rect 17543 33952 18052 33980
rect 17543 33949 17555 33952
rect 17497 33943 17555 33949
rect 18046 33940 18052 33952
rect 18104 33940 18110 33992
rect 11238 33844 11244 33856
rect 11199 33816 11244 33844
rect 11238 33804 11244 33816
rect 11296 33804 11302 33856
rect 13538 33844 13544 33856
rect 13499 33816 13544 33844
rect 13538 33804 13544 33816
rect 13596 33804 13602 33856
rect 17954 33804 17960 33856
rect 18012 33844 18018 33856
rect 18524 33844 18552 34088
rect 20714 34076 20720 34088
rect 20772 34076 20778 34128
rect 21910 34076 21916 34128
rect 21968 34076 21974 34128
rect 23566 34008 23572 34060
rect 23624 34048 23630 34060
rect 23661 34051 23719 34057
rect 23661 34048 23673 34051
rect 23624 34020 23673 34048
rect 23624 34008 23630 34020
rect 23661 34017 23673 34020
rect 23707 34017 23719 34051
rect 23661 34011 23719 34017
rect 20990 33980 20996 33992
rect 20951 33952 20996 33980
rect 20990 33940 20996 33952
rect 21048 33940 21054 33992
rect 21361 33983 21419 33989
rect 21361 33949 21373 33983
rect 21407 33980 21419 33983
rect 21634 33980 21640 33992
rect 21407 33952 21640 33980
rect 21407 33949 21419 33952
rect 21361 33943 21419 33949
rect 21634 33940 21640 33952
rect 21692 33940 21698 33992
rect 23934 33980 23940 33992
rect 23895 33952 23940 33980
rect 23934 33940 23940 33952
rect 23992 33940 23998 33992
rect 18012 33816 18552 33844
rect 18923 33847 18981 33853
rect 18012 33804 18018 33816
rect 18923 33813 18935 33847
rect 18969 33844 18981 33847
rect 19334 33844 19340 33856
rect 18969 33816 19340 33844
rect 18969 33813 18981 33816
rect 18923 33807 18981 33813
rect 19334 33804 19340 33816
rect 19392 33804 19398 33856
rect 21174 33804 21180 33856
rect 21232 33844 21238 33856
rect 22787 33847 22845 33853
rect 22787 33844 22799 33847
rect 21232 33816 22799 33844
rect 21232 33804 21238 33816
rect 22787 33813 22799 33816
rect 22833 33844 22845 33847
rect 23566 33844 23572 33856
rect 22833 33816 23572 33844
rect 22833 33813 22845 33816
rect 22787 33807 22845 33813
rect 23566 33804 23572 33816
rect 23624 33804 23630 33856
rect 1104 33754 34316 33776
rect 1104 33702 6517 33754
rect 6569 33702 6581 33754
rect 6633 33702 6645 33754
rect 6697 33702 6709 33754
rect 6761 33702 17588 33754
rect 17640 33702 17652 33754
rect 17704 33702 17716 33754
rect 17768 33702 17780 33754
rect 17832 33702 28658 33754
rect 28710 33702 28722 33754
rect 28774 33702 28786 33754
rect 28838 33702 28850 33754
rect 28902 33702 34316 33754
rect 1104 33680 34316 33702
rect 8202 33640 8208 33652
rect 8163 33612 8208 33640
rect 8202 33600 8208 33612
rect 8260 33600 8266 33652
rect 12526 33600 12532 33652
rect 12584 33640 12590 33652
rect 12805 33643 12863 33649
rect 12805 33640 12817 33643
rect 12584 33612 12817 33640
rect 12584 33600 12590 33612
rect 12805 33609 12817 33612
rect 12851 33609 12863 33643
rect 12805 33603 12863 33609
rect 18046 33600 18052 33652
rect 18104 33640 18110 33652
rect 18141 33643 18199 33649
rect 18141 33640 18153 33643
rect 18104 33612 18153 33640
rect 18104 33600 18110 33612
rect 18141 33609 18153 33612
rect 18187 33609 18199 33643
rect 19426 33640 19432 33652
rect 19387 33612 19432 33640
rect 18141 33603 18199 33609
rect 19426 33600 19432 33612
rect 19484 33600 19490 33652
rect 21634 33640 21640 33652
rect 21595 33612 21640 33640
rect 21634 33600 21640 33612
rect 21692 33600 21698 33652
rect 16117 33575 16175 33581
rect 16117 33541 16129 33575
rect 16163 33572 16175 33575
rect 21818 33572 21824 33584
rect 16163 33544 21824 33572
rect 16163 33541 16175 33544
rect 16117 33535 16175 33541
rect 21818 33532 21824 33544
rect 21876 33532 21882 33584
rect 3881 33507 3939 33513
rect 3881 33473 3893 33507
rect 3927 33504 3939 33507
rect 5074 33504 5080 33516
rect 3927 33476 5080 33504
rect 3927 33473 3939 33476
rect 3881 33467 3939 33473
rect 5074 33464 5080 33476
rect 5132 33464 5138 33516
rect 7653 33507 7711 33513
rect 7653 33473 7665 33507
rect 7699 33504 7711 33507
rect 12161 33507 12219 33513
rect 12161 33504 12173 33507
rect 7699 33476 12173 33504
rect 7699 33473 7711 33476
rect 7653 33467 7711 33473
rect 12161 33473 12173 33476
rect 12207 33473 12219 33507
rect 12161 33467 12219 33473
rect 12345 33507 12403 33513
rect 12345 33473 12357 33507
rect 12391 33504 12403 33507
rect 13538 33504 13544 33516
rect 12391 33476 13544 33504
rect 12391 33473 12403 33476
rect 12345 33467 12403 33473
rect 2958 33396 2964 33448
rect 3016 33436 3022 33448
rect 3697 33439 3755 33445
rect 3697 33436 3709 33439
rect 3016 33408 3709 33436
rect 3016 33396 3022 33408
rect 3697 33405 3709 33408
rect 3743 33405 3755 33439
rect 3697 33399 3755 33405
rect 3789 33439 3847 33445
rect 3789 33405 3801 33439
rect 3835 33405 3847 33439
rect 3970 33436 3976 33448
rect 3931 33408 3976 33436
rect 3789 33399 3847 33405
rect 3050 33328 3056 33380
rect 3108 33368 3114 33380
rect 3804 33368 3832 33399
rect 3970 33396 3976 33408
rect 4028 33396 4034 33448
rect 8662 33436 8668 33448
rect 8623 33408 8668 33436
rect 8662 33396 8668 33408
rect 8720 33396 8726 33448
rect 8938 33436 8944 33448
rect 8899 33408 8944 33436
rect 8938 33396 8944 33408
rect 8996 33396 9002 33448
rect 9490 33436 9496 33448
rect 9451 33408 9496 33436
rect 9490 33396 9496 33408
rect 9548 33396 9554 33448
rect 10410 33396 10416 33448
rect 10468 33436 10474 33448
rect 10505 33439 10563 33445
rect 10505 33436 10517 33439
rect 10468 33408 10517 33436
rect 10468 33396 10474 33408
rect 10505 33405 10517 33408
rect 10551 33405 10563 33439
rect 12176 33436 12204 33467
rect 13538 33464 13544 33476
rect 13596 33464 13602 33516
rect 13814 33464 13820 33516
rect 13872 33504 13878 33516
rect 14369 33507 14427 33513
rect 14369 33504 14381 33507
rect 13872 33476 14381 33504
rect 13872 33464 13878 33476
rect 14369 33473 14381 33476
rect 14415 33473 14427 33507
rect 14369 33467 14427 33473
rect 18785 33507 18843 33513
rect 18785 33473 18797 33507
rect 18831 33473 18843 33507
rect 19886 33504 19892 33516
rect 19847 33476 19892 33504
rect 18785 33467 18843 33473
rect 12526 33436 12532 33448
rect 12176 33408 12532 33436
rect 10505 33399 10563 33405
rect 12526 33396 12532 33408
rect 12584 33396 12590 33448
rect 13262 33436 13268 33448
rect 13223 33408 13268 33436
rect 13262 33396 13268 33408
rect 13320 33396 13326 33448
rect 13446 33436 13452 33448
rect 13359 33408 13452 33436
rect 13446 33396 13452 33408
rect 13504 33396 13510 33448
rect 18598 33396 18604 33448
rect 18656 33436 18662 33448
rect 18800 33436 18828 33467
rect 19886 33464 19892 33476
rect 19944 33464 19950 33516
rect 20073 33507 20131 33513
rect 20073 33473 20085 33507
rect 20119 33504 20131 33507
rect 20714 33504 20720 33516
rect 20119 33476 20720 33504
rect 20119 33473 20131 33476
rect 20073 33467 20131 33473
rect 20088 33436 20116 33467
rect 20714 33464 20720 33476
rect 20772 33504 20778 33516
rect 20993 33507 21051 33513
rect 20993 33504 21005 33507
rect 20772 33476 21005 33504
rect 20772 33464 20778 33476
rect 20993 33473 21005 33476
rect 21039 33473 21051 33507
rect 21174 33504 21180 33516
rect 21135 33476 21180 33504
rect 20993 33467 21051 33473
rect 21174 33464 21180 33476
rect 21232 33464 21238 33516
rect 25314 33436 25320 33448
rect 18656 33408 20116 33436
rect 25275 33408 25320 33436
rect 18656 33396 18662 33408
rect 25314 33396 25320 33408
rect 25372 33396 25378 33448
rect 25685 33439 25743 33445
rect 25685 33405 25697 33439
rect 25731 33436 25743 33439
rect 27798 33436 27804 33448
rect 25731 33408 27804 33436
rect 25731 33405 25743 33408
rect 25685 33399 25743 33405
rect 27798 33396 27804 33408
rect 27856 33436 27862 33448
rect 27893 33439 27951 33445
rect 27893 33436 27905 33439
rect 27856 33408 27905 33436
rect 27856 33396 27862 33408
rect 27893 33405 27905 33408
rect 27939 33405 27951 33439
rect 27893 33399 27951 33405
rect 29270 33396 29276 33448
rect 29328 33396 29334 33448
rect 33594 33436 33600 33448
rect 33555 33408 33600 33436
rect 33594 33396 33600 33408
rect 33652 33396 33658 33448
rect 5442 33368 5448 33380
rect 3108 33340 5448 33368
rect 3108 33328 3114 33340
rect 5442 33328 5448 33340
rect 5500 33328 5506 33380
rect 9950 33328 9956 33380
rect 10008 33368 10014 33380
rect 10321 33371 10379 33377
rect 10321 33368 10333 33371
rect 10008 33340 10333 33368
rect 10008 33328 10014 33340
rect 10321 33337 10333 33340
rect 10367 33337 10379 33371
rect 10321 33331 10379 33337
rect 12437 33371 12495 33377
rect 12437 33337 12449 33371
rect 12483 33368 12495 33371
rect 13357 33371 13415 33377
rect 13357 33368 13369 33371
rect 12483 33340 13369 33368
rect 12483 33337 12495 33340
rect 12437 33331 12495 33337
rect 13357 33337 13369 33340
rect 13403 33337 13415 33371
rect 13357 33331 13415 33337
rect 3513 33303 3571 33309
rect 3513 33269 3525 33303
rect 3559 33300 3571 33303
rect 3602 33300 3608 33312
rect 3559 33272 3608 33300
rect 3559 33269 3571 33272
rect 3513 33263 3571 33269
rect 3602 33260 3608 33272
rect 3660 33260 3666 33312
rect 6914 33260 6920 33312
rect 6972 33300 6978 33312
rect 7742 33300 7748 33312
rect 6972 33272 7748 33300
rect 6972 33260 6978 33272
rect 7742 33260 7748 33272
rect 7800 33260 7806 33312
rect 7837 33303 7895 33309
rect 7837 33269 7849 33303
rect 7883 33300 7895 33303
rect 8570 33300 8576 33312
rect 7883 33272 8576 33300
rect 7883 33269 7895 33272
rect 7837 33263 7895 33269
rect 8570 33260 8576 33272
rect 8628 33260 8634 33312
rect 8754 33300 8760 33312
rect 8715 33272 8760 33300
rect 8754 33260 8760 33272
rect 8812 33260 8818 33312
rect 11238 33260 11244 33312
rect 11296 33300 11302 33312
rect 13464 33300 13492 33396
rect 14645 33371 14703 33377
rect 14645 33337 14657 33371
rect 14691 33368 14703 33371
rect 14734 33368 14740 33380
rect 14691 33340 14740 33368
rect 14691 33337 14703 33340
rect 14645 33331 14703 33337
rect 14734 33328 14740 33340
rect 14792 33328 14798 33380
rect 15488 33312 15516 33354
rect 21910 33328 21916 33380
rect 21968 33368 21974 33380
rect 24302 33368 24308 33380
rect 21968 33340 24308 33368
rect 21968 33328 21974 33340
rect 24302 33328 24308 33340
rect 24360 33328 24366 33380
rect 28166 33368 28172 33380
rect 28127 33340 28172 33368
rect 28166 33328 28172 33340
rect 28224 33328 28230 33380
rect 29917 33371 29975 33377
rect 29917 33337 29929 33371
rect 29963 33368 29975 33371
rect 30006 33368 30012 33380
rect 29963 33340 30012 33368
rect 29963 33337 29975 33340
rect 29917 33331 29975 33337
rect 30006 33328 30012 33340
rect 30064 33328 30070 33380
rect 11296 33272 13492 33300
rect 11296 33260 11302 33272
rect 15470 33260 15476 33312
rect 15528 33260 15534 33312
rect 18506 33300 18512 33312
rect 18467 33272 18512 33300
rect 18506 33260 18512 33272
rect 18564 33260 18570 33312
rect 18601 33303 18659 33309
rect 18601 33269 18613 33303
rect 18647 33300 18659 33303
rect 19334 33300 19340 33312
rect 18647 33272 19340 33300
rect 18647 33269 18659 33272
rect 18601 33263 18659 33269
rect 19334 33260 19340 33272
rect 19392 33300 19398 33312
rect 19794 33300 19800 33312
rect 19392 33272 19800 33300
rect 19392 33260 19398 33272
rect 19794 33260 19800 33272
rect 19852 33260 19858 33312
rect 21266 33300 21272 33312
rect 21227 33272 21272 33300
rect 21266 33260 21272 33272
rect 21324 33260 21330 33312
rect 23658 33260 23664 33312
rect 23716 33300 23722 33312
rect 23891 33303 23949 33309
rect 23891 33300 23903 33303
rect 23716 33272 23903 33300
rect 23716 33260 23722 33272
rect 23891 33269 23903 33272
rect 23937 33269 23949 33303
rect 33410 33300 33416 33312
rect 33371 33272 33416 33300
rect 23891 33263 23949 33269
rect 33410 33260 33416 33272
rect 33468 33260 33474 33312
rect 1104 33210 34316 33232
rect 1104 33158 12052 33210
rect 12104 33158 12116 33210
rect 12168 33158 12180 33210
rect 12232 33158 12244 33210
rect 12296 33158 23123 33210
rect 23175 33158 23187 33210
rect 23239 33158 23251 33210
rect 23303 33158 23315 33210
rect 23367 33158 34316 33210
rect 1104 33136 34316 33158
rect 1581 33099 1639 33105
rect 1581 33065 1593 33099
rect 1627 33096 1639 33099
rect 7650 33096 7656 33108
rect 1627 33068 7656 33096
rect 1627 33065 1639 33068
rect 1581 33059 1639 33065
rect 7650 33056 7656 33068
rect 7708 33056 7714 33108
rect 7742 33056 7748 33108
rect 7800 33056 7806 33108
rect 10502 33096 10508 33108
rect 10463 33068 10508 33096
rect 10502 33056 10508 33068
rect 10560 33056 10566 33108
rect 12437 33099 12495 33105
rect 12437 33065 12449 33099
rect 12483 33065 12495 33099
rect 12437 33059 12495 33065
rect 3878 32988 3884 33040
rect 3936 33028 3942 33040
rect 7760 33028 7788 33056
rect 12452 33028 12480 33059
rect 17402 33056 17408 33108
rect 17460 33096 17466 33108
rect 17460 33068 17816 33096
rect 17460 33056 17466 33068
rect 17788 33040 17816 33068
rect 3936 33000 6914 33028
rect 7760 33000 8432 33028
rect 3936 32988 3942 33000
rect 1394 32960 1400 32972
rect 1355 32932 1400 32960
rect 1394 32920 1400 32932
rect 1452 32920 1458 32972
rect 5626 32960 5632 32972
rect 5684 32969 5690 32972
rect 5920 32969 5948 33000
rect 5596 32932 5632 32960
rect 5626 32920 5632 32932
rect 5684 32923 5696 32969
rect 5905 32963 5963 32969
rect 5905 32929 5917 32963
rect 5951 32929 5963 32963
rect 5905 32923 5963 32929
rect 5684 32920 5690 32923
rect 6886 32824 6914 33000
rect 7673 32963 7731 32969
rect 7673 32929 7685 32963
rect 7719 32960 7731 32963
rect 8294 32960 8300 32972
rect 7719 32932 8300 32960
rect 7719 32929 7731 32932
rect 7673 32923 7731 32929
rect 8294 32920 8300 32932
rect 8352 32920 8358 32972
rect 8404 32969 8432 33000
rect 9600 33000 12480 33028
rect 9600 32969 9628 33000
rect 17770 32988 17776 33040
rect 17828 32988 17834 33040
rect 18187 33031 18245 33037
rect 18187 32997 18199 33031
rect 18233 33028 18245 33031
rect 18506 33028 18512 33040
rect 18233 33000 18512 33028
rect 18233 32997 18245 33000
rect 18187 32991 18245 32997
rect 18506 32988 18512 33000
rect 18564 33028 18570 33040
rect 19981 33031 20039 33037
rect 19981 33028 19993 33031
rect 18564 33000 19993 33028
rect 18564 32988 18570 33000
rect 19981 32997 19993 33000
rect 20027 32997 20039 33031
rect 23566 33028 23572 33040
rect 23527 33000 23572 33028
rect 19981 32991 20039 32997
rect 23566 32988 23572 33000
rect 23624 32988 23630 33040
rect 8389 32963 8447 32969
rect 8389 32929 8401 32963
rect 8435 32929 8447 32963
rect 8389 32923 8447 32929
rect 9585 32963 9643 32969
rect 9585 32929 9597 32963
rect 9631 32929 9643 32963
rect 9585 32923 9643 32929
rect 10045 32963 10103 32969
rect 10045 32929 10057 32963
rect 10091 32960 10103 32963
rect 10226 32960 10232 32972
rect 10091 32932 10232 32960
rect 10091 32929 10103 32932
rect 10045 32923 10103 32929
rect 10226 32920 10232 32932
rect 10284 32920 10290 32972
rect 10410 32920 10416 32972
rect 10468 32960 10474 32972
rect 10505 32963 10563 32969
rect 10505 32960 10517 32963
rect 10468 32932 10517 32960
rect 10468 32920 10474 32932
rect 10505 32929 10517 32932
rect 10551 32929 10563 32963
rect 10505 32923 10563 32929
rect 10689 32963 10747 32969
rect 10689 32929 10701 32963
rect 10735 32960 10747 32963
rect 11238 32960 11244 32972
rect 10735 32932 11244 32960
rect 10735 32929 10747 32932
rect 10689 32923 10747 32929
rect 7929 32895 7987 32901
rect 7929 32861 7941 32895
rect 7975 32892 7987 32895
rect 9674 32892 9680 32904
rect 7975 32864 9680 32892
rect 7975 32861 7987 32864
rect 7929 32855 7987 32861
rect 6886 32796 7052 32824
rect 4522 32756 4528 32768
rect 4483 32728 4528 32756
rect 4522 32716 4528 32728
rect 4580 32716 4586 32768
rect 6549 32759 6607 32765
rect 6549 32725 6561 32759
rect 6595 32756 6607 32759
rect 6914 32756 6920 32768
rect 6595 32728 6920 32756
rect 6595 32725 6607 32728
rect 6549 32719 6607 32725
rect 6914 32716 6920 32728
rect 6972 32716 6978 32768
rect 7024 32756 7052 32796
rect 7944 32756 7972 32855
rect 9674 32852 9680 32864
rect 9732 32852 9738 32904
rect 9861 32895 9919 32901
rect 9861 32861 9873 32895
rect 9907 32892 9919 32895
rect 9950 32892 9956 32904
rect 9907 32864 9956 32892
rect 9907 32861 9919 32864
rect 9861 32855 9919 32861
rect 9950 32852 9956 32864
rect 10008 32852 10014 32904
rect 10318 32852 10324 32904
rect 10376 32892 10382 32904
rect 10704 32892 10732 32923
rect 11238 32920 11244 32932
rect 11296 32920 11302 32972
rect 12805 32963 12863 32969
rect 12805 32929 12817 32963
rect 12851 32960 12863 32963
rect 13538 32960 13544 32972
rect 12851 32932 13544 32960
rect 12851 32929 12863 32932
rect 12805 32923 12863 32929
rect 13538 32920 13544 32932
rect 13596 32920 13602 32972
rect 14826 32920 14832 32972
rect 14884 32960 14890 32972
rect 15105 32963 15163 32969
rect 15105 32960 15117 32963
rect 14884 32932 15117 32960
rect 14884 32920 14890 32932
rect 15105 32929 15117 32932
rect 15151 32929 15163 32963
rect 15105 32923 15163 32929
rect 16298 32920 16304 32972
rect 16356 32960 16362 32972
rect 16393 32963 16451 32969
rect 16393 32960 16405 32963
rect 16356 32932 16405 32960
rect 16356 32920 16362 32932
rect 16393 32929 16405 32932
rect 16439 32929 16451 32963
rect 16393 32923 16451 32929
rect 23422 32963 23480 32969
rect 23422 32929 23434 32963
rect 23468 32960 23480 32963
rect 23750 32960 23756 32972
rect 23468 32932 23756 32960
rect 23468 32929 23480 32932
rect 23422 32923 23480 32929
rect 23750 32920 23756 32932
rect 23808 32920 23814 32972
rect 33410 32960 33416 32972
rect 33371 32932 33416 32960
rect 33410 32920 33416 32932
rect 33468 32920 33474 32972
rect 12894 32892 12900 32904
rect 10376 32864 10732 32892
rect 12855 32864 12900 32892
rect 10376 32852 10382 32864
rect 12894 32852 12900 32864
rect 12952 32852 12958 32904
rect 12986 32852 12992 32904
rect 13044 32892 13050 32904
rect 15194 32892 15200 32904
rect 13044 32864 13089 32892
rect 15155 32864 15200 32892
rect 13044 32852 13050 32864
rect 15194 32852 15200 32864
rect 15252 32852 15258 32904
rect 15289 32895 15347 32901
rect 15289 32861 15301 32895
rect 15335 32861 15347 32895
rect 15289 32855 15347 32861
rect 16761 32895 16819 32901
rect 16761 32861 16773 32895
rect 16807 32892 16819 32895
rect 17954 32892 17960 32904
rect 16807 32864 17960 32892
rect 16807 32861 16819 32864
rect 16761 32855 16819 32861
rect 13004 32824 13032 32852
rect 15304 32824 15332 32855
rect 17954 32852 17960 32864
rect 18012 32852 18018 32904
rect 19794 32852 19800 32904
rect 19852 32892 19858 32904
rect 20128 32895 20186 32901
rect 20128 32892 20140 32895
rect 19852 32864 20140 32892
rect 19852 32852 19858 32864
rect 20128 32861 20140 32864
rect 20174 32861 20186 32895
rect 20128 32855 20186 32861
rect 20349 32895 20407 32901
rect 20349 32861 20361 32895
rect 20395 32892 20407 32895
rect 21266 32892 21272 32904
rect 20395 32864 21272 32892
rect 20395 32861 20407 32864
rect 20349 32855 20407 32861
rect 21266 32852 21272 32864
rect 21324 32852 21330 32904
rect 22830 32852 22836 32904
rect 22888 32892 22894 32904
rect 23201 32895 23259 32901
rect 23201 32892 23213 32895
rect 22888 32864 23213 32892
rect 22888 32852 22894 32864
rect 23201 32861 23213 32864
rect 23247 32861 23259 32895
rect 23201 32855 23259 32861
rect 13004 32796 15332 32824
rect 19150 32784 19156 32836
rect 19208 32824 19214 32836
rect 22925 32827 22983 32833
rect 22925 32824 22937 32827
rect 19208 32796 22937 32824
rect 19208 32784 19214 32796
rect 22925 32793 22937 32796
rect 22971 32793 22983 32827
rect 22925 32787 22983 32793
rect 23293 32827 23351 32833
rect 23293 32793 23305 32827
rect 23339 32824 23351 32827
rect 23658 32824 23664 32836
rect 23339 32796 23664 32824
rect 23339 32793 23351 32796
rect 23293 32787 23351 32793
rect 23658 32784 23664 32796
rect 23716 32784 23722 32836
rect 8478 32756 8484 32768
rect 7024 32728 7972 32756
rect 8439 32728 8484 32756
rect 8478 32716 8484 32728
rect 8536 32716 8542 32768
rect 8938 32716 8944 32768
rect 8996 32756 9002 32768
rect 9582 32756 9588 32768
rect 8996 32728 9588 32756
rect 8996 32716 9002 32728
rect 9582 32716 9588 32728
rect 9640 32756 9646 32768
rect 9723 32759 9781 32765
rect 9723 32756 9735 32759
rect 9640 32728 9735 32756
rect 9640 32716 9646 32728
rect 9723 32725 9735 32728
rect 9769 32725 9781 32759
rect 9723 32719 9781 32725
rect 9953 32759 10011 32765
rect 9953 32725 9965 32759
rect 9999 32756 10011 32759
rect 10042 32756 10048 32768
rect 9999 32728 10048 32756
rect 9999 32725 10011 32728
rect 9953 32719 10011 32725
rect 10042 32716 10048 32728
rect 10100 32716 10106 32768
rect 14182 32716 14188 32768
rect 14240 32756 14246 32768
rect 14737 32759 14795 32765
rect 14737 32756 14749 32759
rect 14240 32728 14749 32756
rect 14240 32716 14246 32728
rect 14737 32725 14749 32728
rect 14783 32725 14795 32759
rect 14737 32719 14795 32725
rect 19886 32716 19892 32768
rect 19944 32756 19950 32768
rect 20254 32756 20260 32768
rect 19944 32728 20260 32756
rect 19944 32716 19950 32728
rect 20254 32716 20260 32728
rect 20312 32716 20318 32768
rect 20438 32756 20444 32768
rect 20399 32728 20444 32756
rect 20438 32716 20444 32728
rect 20496 32716 20502 32768
rect 33502 32756 33508 32768
rect 33463 32728 33508 32756
rect 33502 32716 33508 32728
rect 33560 32716 33566 32768
rect 1104 32666 34316 32688
rect 1104 32614 6517 32666
rect 6569 32614 6581 32666
rect 6633 32614 6645 32666
rect 6697 32614 6709 32666
rect 6761 32614 17588 32666
rect 17640 32614 17652 32666
rect 17704 32614 17716 32666
rect 17768 32614 17780 32666
rect 17832 32614 28658 32666
rect 28710 32614 28722 32666
rect 28774 32614 28786 32666
rect 28838 32614 28850 32666
rect 28902 32614 34316 32666
rect 1104 32592 34316 32614
rect 5074 32552 5080 32564
rect 5035 32524 5080 32552
rect 5074 32512 5080 32524
rect 5132 32512 5138 32564
rect 8294 32552 8300 32564
rect 8255 32524 8300 32552
rect 8294 32512 8300 32524
rect 8352 32512 8358 32564
rect 8570 32512 8576 32564
rect 8628 32552 8634 32564
rect 9033 32555 9091 32561
rect 9033 32552 9045 32555
rect 8628 32524 9045 32552
rect 8628 32512 8634 32524
rect 9033 32521 9045 32524
rect 9079 32521 9091 32555
rect 9033 32515 9091 32521
rect 12894 32512 12900 32564
rect 12952 32552 12958 32564
rect 13081 32555 13139 32561
rect 13081 32552 13093 32555
rect 12952 32524 13093 32552
rect 12952 32512 12958 32524
rect 13081 32521 13093 32524
rect 13127 32521 13139 32555
rect 13538 32552 13544 32564
rect 13499 32524 13544 32552
rect 13081 32515 13139 32521
rect 5350 32376 5356 32428
rect 5408 32416 5414 32428
rect 5721 32419 5779 32425
rect 5721 32416 5733 32419
rect 5408 32388 5733 32416
rect 5408 32376 5414 32388
rect 5721 32385 5733 32388
rect 5767 32416 5779 32419
rect 7466 32416 7472 32428
rect 5767 32388 7472 32416
rect 5767 32385 5779 32388
rect 5721 32379 5779 32385
rect 7466 32376 7472 32388
rect 7524 32376 7530 32428
rect 12526 32416 12532 32428
rect 8496 32388 9076 32416
rect 12487 32388 12532 32416
rect 8496 32360 8524 32388
rect 3602 32308 3608 32360
rect 3660 32357 3666 32360
rect 3660 32348 3672 32357
rect 3878 32348 3884 32360
rect 3660 32320 3705 32348
rect 3839 32320 3884 32348
rect 3660 32311 3672 32320
rect 3660 32308 3666 32311
rect 3878 32308 3884 32320
rect 3936 32308 3942 32360
rect 5445 32351 5503 32357
rect 5445 32317 5457 32351
rect 5491 32348 5503 32351
rect 6914 32348 6920 32360
rect 5491 32320 6920 32348
rect 5491 32317 5503 32320
rect 5445 32311 5503 32317
rect 6914 32308 6920 32320
rect 6972 32308 6978 32360
rect 8478 32348 8484 32360
rect 8439 32320 8484 32348
rect 8478 32308 8484 32320
rect 8536 32308 8542 32360
rect 9048 32357 9076 32388
rect 12526 32376 12532 32388
rect 12584 32376 12590 32428
rect 8573 32351 8631 32357
rect 8573 32317 8585 32351
rect 8619 32348 8631 32351
rect 9033 32351 9091 32357
rect 8619 32320 8984 32348
rect 8619 32317 8631 32320
rect 8573 32311 8631 32317
rect 8297 32283 8355 32289
rect 8297 32249 8309 32283
rect 8343 32280 8355 32283
rect 8754 32280 8760 32292
rect 8343 32252 8760 32280
rect 8343 32249 8355 32252
rect 8297 32243 8355 32249
rect 8754 32240 8760 32252
rect 8812 32240 8818 32292
rect 8956 32280 8984 32320
rect 9033 32317 9045 32351
rect 9079 32317 9091 32351
rect 9033 32311 9091 32317
rect 9217 32351 9275 32357
rect 9217 32317 9229 32351
rect 9263 32348 9275 32351
rect 9582 32348 9588 32360
rect 9263 32320 9588 32348
rect 9263 32317 9275 32320
rect 9217 32311 9275 32317
rect 9582 32308 9588 32320
rect 9640 32308 9646 32360
rect 9674 32308 9680 32360
rect 9732 32348 9738 32360
rect 10042 32357 10048 32360
rect 9769 32351 9827 32357
rect 9769 32348 9781 32351
rect 9732 32320 9781 32348
rect 9732 32308 9738 32320
rect 9769 32317 9781 32320
rect 9815 32317 9827 32351
rect 10036 32348 10048 32357
rect 10003 32320 10048 32348
rect 9769 32311 9827 32317
rect 10036 32311 10048 32320
rect 10042 32308 10048 32311
rect 10100 32308 10106 32360
rect 13096 32348 13124 32515
rect 13538 32512 13544 32524
rect 13596 32512 13602 32564
rect 14826 32552 14832 32564
rect 14787 32524 14832 32552
rect 14826 32512 14832 32524
rect 14884 32512 14890 32564
rect 33502 32552 33508 32564
rect 16546 32524 33508 32552
rect 16546 32484 16574 32524
rect 33502 32512 33508 32524
rect 33560 32512 33566 32564
rect 17954 32484 17960 32496
rect 14016 32456 16574 32484
rect 17915 32456 17960 32484
rect 14016 32425 14044 32456
rect 17954 32444 17960 32456
rect 18012 32444 18018 32496
rect 19334 32484 19340 32496
rect 19295 32456 19340 32484
rect 19334 32444 19340 32456
rect 19392 32444 19398 32496
rect 21266 32444 21272 32496
rect 21324 32484 21330 32496
rect 21591 32487 21649 32493
rect 21591 32484 21603 32487
rect 21324 32456 21603 32484
rect 21324 32444 21330 32456
rect 21591 32453 21603 32456
rect 21637 32453 21649 32487
rect 21591 32447 21649 32453
rect 24765 32487 24823 32493
rect 24765 32453 24777 32487
rect 24811 32484 24823 32487
rect 25314 32484 25320 32496
rect 24811 32456 25320 32484
rect 24811 32453 24823 32456
rect 24765 32447 24823 32453
rect 25314 32444 25320 32456
rect 25372 32444 25378 32496
rect 28166 32444 28172 32496
rect 28224 32484 28230 32496
rect 28905 32487 28963 32493
rect 28905 32484 28917 32487
rect 28224 32456 28917 32484
rect 28224 32444 28230 32456
rect 28905 32453 28917 32456
rect 28951 32453 28963 32487
rect 28905 32447 28963 32453
rect 14001 32419 14059 32425
rect 14001 32385 14013 32419
rect 14047 32385 14059 32419
rect 14001 32379 14059 32385
rect 14093 32419 14151 32425
rect 14093 32385 14105 32419
rect 14139 32385 14151 32419
rect 15286 32416 15292 32428
rect 15247 32388 15292 32416
rect 14093 32379 14151 32385
rect 13909 32351 13967 32357
rect 13909 32348 13921 32351
rect 13096 32320 13921 32348
rect 13909 32317 13921 32320
rect 13955 32317 13967 32351
rect 14108 32348 14136 32379
rect 15286 32376 15292 32388
rect 15344 32376 15350 32428
rect 15381 32419 15439 32425
rect 15381 32385 15393 32419
rect 15427 32385 15439 32419
rect 15381 32379 15439 32385
rect 15194 32348 15200 32360
rect 13909 32311 13967 32317
rect 14016 32320 14136 32348
rect 15155 32320 15200 32348
rect 9950 32280 9956 32292
rect 8956 32252 9956 32280
rect 9950 32240 9956 32252
rect 10008 32240 10014 32292
rect 13262 32280 13268 32292
rect 10060 32252 13268 32280
rect 2501 32215 2559 32221
rect 2501 32181 2513 32215
rect 2547 32212 2559 32215
rect 3142 32212 3148 32224
rect 2547 32184 3148 32212
rect 2547 32181 2559 32184
rect 2501 32175 2559 32181
rect 3142 32172 3148 32184
rect 3200 32172 3206 32224
rect 4522 32172 4528 32224
rect 4580 32212 4586 32224
rect 5534 32212 5540 32224
rect 4580 32184 5540 32212
rect 4580 32172 4586 32184
rect 5534 32172 5540 32184
rect 5592 32172 5598 32224
rect 5718 32172 5724 32224
rect 5776 32212 5782 32224
rect 6917 32215 6975 32221
rect 6917 32212 6929 32215
rect 5776 32184 6929 32212
rect 5776 32172 5782 32184
rect 6917 32181 6929 32184
rect 6963 32181 6975 32215
rect 7282 32212 7288 32224
rect 7243 32184 7288 32212
rect 6917 32175 6975 32181
rect 7282 32172 7288 32184
rect 7340 32172 7346 32224
rect 7374 32172 7380 32224
rect 7432 32212 7438 32224
rect 7432 32184 7477 32212
rect 7432 32172 7438 32184
rect 9582 32172 9588 32224
rect 9640 32212 9646 32224
rect 10060 32212 10088 32252
rect 13262 32240 13268 32252
rect 13320 32240 13326 32292
rect 14016 32280 14044 32320
rect 15194 32308 15200 32320
rect 15252 32308 15258 32360
rect 15396 32348 15424 32379
rect 18138 32376 18144 32428
rect 18196 32416 18202 32428
rect 18598 32416 18604 32428
rect 18196 32388 18604 32416
rect 18196 32376 18202 32388
rect 18598 32376 18604 32388
rect 18656 32376 18662 32428
rect 20438 32416 20444 32428
rect 19352 32388 20444 32416
rect 19150 32348 19156 32360
rect 15304 32320 15424 32348
rect 19111 32320 19156 32348
rect 15304 32280 15332 32320
rect 19150 32308 19156 32320
rect 19208 32308 19214 32360
rect 19352 32357 19380 32388
rect 20438 32376 20444 32388
rect 20496 32376 20502 32428
rect 22741 32419 22799 32425
rect 22741 32385 22753 32419
rect 22787 32416 22799 32419
rect 23474 32416 23480 32428
rect 22787 32388 23480 32416
rect 22787 32385 22799 32388
rect 22741 32379 22799 32385
rect 23474 32376 23480 32388
rect 23532 32416 23538 32428
rect 23934 32416 23940 32428
rect 23532 32388 23940 32416
rect 23532 32376 23538 32388
rect 23934 32376 23940 32388
rect 23992 32416 23998 32428
rect 24213 32419 24271 32425
rect 24213 32416 24225 32419
rect 23992 32388 24225 32416
rect 23992 32376 23998 32388
rect 24213 32385 24225 32388
rect 24259 32416 24271 32419
rect 26513 32419 26571 32425
rect 26513 32416 26525 32419
rect 24259 32388 26525 32416
rect 24259 32385 24271 32388
rect 24213 32379 24271 32385
rect 26513 32385 26525 32388
rect 26559 32416 26571 32419
rect 26602 32416 26608 32428
rect 26559 32388 26608 32416
rect 26559 32385 26571 32388
rect 26513 32379 26571 32385
rect 26602 32376 26608 32388
rect 26660 32376 26666 32428
rect 29454 32416 29460 32428
rect 29415 32388 29460 32416
rect 29454 32376 29460 32388
rect 29512 32376 29518 32428
rect 19337 32351 19395 32357
rect 19337 32317 19349 32351
rect 19383 32317 19395 32351
rect 19337 32311 19395 32317
rect 19797 32351 19855 32357
rect 19797 32317 19809 32351
rect 19843 32317 19855 32351
rect 20162 32348 20168 32360
rect 20123 32320 20168 32348
rect 19797 32311 19855 32317
rect 14016 32252 15332 32280
rect 18417 32283 18475 32289
rect 11146 32212 11152 32224
rect 9640 32184 10088 32212
rect 11107 32184 11152 32212
rect 9640 32172 9646 32184
rect 11146 32172 11152 32184
rect 11204 32172 11210 32224
rect 12434 32172 12440 32224
rect 12492 32212 12498 32224
rect 12621 32215 12679 32221
rect 12621 32212 12633 32215
rect 12492 32184 12633 32212
rect 12492 32172 12498 32184
rect 12621 32181 12633 32184
rect 12667 32181 12679 32215
rect 12621 32175 12679 32181
rect 12713 32215 12771 32221
rect 12713 32181 12725 32215
rect 12759 32212 12771 32215
rect 12986 32212 12992 32224
rect 12759 32184 12992 32212
rect 12759 32181 12771 32184
rect 12713 32175 12771 32181
rect 12986 32172 12992 32184
rect 13044 32172 13050 32224
rect 13170 32172 13176 32224
rect 13228 32212 13234 32224
rect 14016 32212 14044 32252
rect 18417 32249 18429 32283
rect 18463 32280 18475 32283
rect 18506 32280 18512 32292
rect 18463 32252 18512 32280
rect 18463 32249 18475 32252
rect 18417 32243 18475 32249
rect 18506 32240 18512 32252
rect 18564 32240 18570 32292
rect 13228 32184 14044 32212
rect 13228 32172 13234 32184
rect 17954 32172 17960 32224
rect 18012 32212 18018 32224
rect 18325 32215 18383 32221
rect 18325 32212 18337 32215
rect 18012 32184 18337 32212
rect 18012 32172 18018 32184
rect 18325 32181 18337 32184
rect 18371 32181 18383 32215
rect 19812 32212 19840 32311
rect 20162 32308 20168 32320
rect 20220 32308 20226 32360
rect 22925 32351 22983 32357
rect 22925 32317 22937 32351
rect 22971 32348 22983 32351
rect 23658 32348 23664 32360
rect 22971 32320 23664 32348
rect 22971 32317 22983 32320
rect 22925 32311 22983 32317
rect 23658 32308 23664 32320
rect 23716 32348 23722 32360
rect 24305 32351 24363 32357
rect 24305 32348 24317 32351
rect 23716 32320 24317 32348
rect 23716 32308 23722 32320
rect 24305 32317 24317 32320
rect 24351 32317 24363 32351
rect 24305 32311 24363 32317
rect 27798 32308 27804 32360
rect 27856 32348 27862 32360
rect 30101 32351 30159 32357
rect 30101 32348 30113 32351
rect 27856 32320 30113 32348
rect 27856 32308 27862 32320
rect 30101 32317 30113 32320
rect 30147 32317 30159 32351
rect 30101 32311 30159 32317
rect 21174 32240 21180 32292
rect 21232 32280 21238 32292
rect 21910 32280 21916 32292
rect 21232 32252 21916 32280
rect 21232 32240 21238 32252
rect 21910 32240 21916 32252
rect 21968 32240 21974 32292
rect 23750 32240 23756 32292
rect 23808 32280 23814 32292
rect 24397 32283 24455 32289
rect 24397 32280 24409 32283
rect 23808 32252 24409 32280
rect 23808 32240 23814 32252
rect 24397 32249 24409 32252
rect 24443 32249 24455 32283
rect 24397 32243 24455 32249
rect 26329 32283 26387 32289
rect 26329 32249 26341 32283
rect 26375 32280 26387 32283
rect 26694 32280 26700 32292
rect 26375 32252 26700 32280
rect 26375 32249 26387 32252
rect 26329 32243 26387 32249
rect 26694 32240 26700 32252
rect 26752 32240 26758 32292
rect 30377 32283 30435 32289
rect 30377 32249 30389 32283
rect 30423 32280 30435 32283
rect 30466 32280 30472 32292
rect 30423 32252 30472 32280
rect 30423 32249 30435 32252
rect 30377 32243 30435 32249
rect 30466 32240 30472 32252
rect 30524 32240 30530 32292
rect 30650 32240 30656 32292
rect 30708 32280 30714 32292
rect 30708 32252 30866 32280
rect 30708 32240 30714 32252
rect 20990 32212 20996 32224
rect 19812 32184 20996 32212
rect 18325 32175 18383 32181
rect 20990 32172 20996 32184
rect 21048 32212 21054 32224
rect 21358 32212 21364 32224
rect 21048 32184 21364 32212
rect 21048 32172 21054 32184
rect 21358 32172 21364 32184
rect 21416 32172 21422 32224
rect 22094 32172 22100 32224
rect 22152 32212 22158 32224
rect 22830 32212 22836 32224
rect 22152 32184 22836 32212
rect 22152 32172 22158 32184
rect 22830 32172 22836 32184
rect 22888 32172 22894 32224
rect 23014 32172 23020 32224
rect 23072 32212 23078 32224
rect 23293 32215 23351 32221
rect 23293 32212 23305 32215
rect 23072 32184 23305 32212
rect 23072 32172 23078 32184
rect 23293 32181 23305 32184
rect 23339 32181 23351 32215
rect 25866 32212 25872 32224
rect 25827 32184 25872 32212
rect 23293 32175 23351 32181
rect 25866 32172 25872 32184
rect 25924 32172 25930 32224
rect 26234 32172 26240 32224
rect 26292 32212 26298 32224
rect 29270 32212 29276 32224
rect 26292 32184 26337 32212
rect 29231 32184 29276 32212
rect 26292 32172 26298 32184
rect 29270 32172 29276 32184
rect 29328 32172 29334 32224
rect 29365 32215 29423 32221
rect 29365 32181 29377 32215
rect 29411 32212 29423 32215
rect 30742 32212 30748 32224
rect 29411 32184 30748 32212
rect 29411 32181 29423 32184
rect 29365 32175 29423 32181
rect 30742 32172 30748 32184
rect 30800 32212 30806 32224
rect 31849 32215 31907 32221
rect 31849 32212 31861 32215
rect 30800 32184 31861 32212
rect 30800 32172 30806 32184
rect 31849 32181 31861 32184
rect 31895 32181 31907 32215
rect 31849 32175 31907 32181
rect 1104 32122 34316 32144
rect 1104 32070 12052 32122
rect 12104 32070 12116 32122
rect 12168 32070 12180 32122
rect 12232 32070 12244 32122
rect 12296 32070 23123 32122
rect 23175 32070 23187 32122
rect 23239 32070 23251 32122
rect 23303 32070 23315 32122
rect 23367 32070 34316 32122
rect 1104 32048 34316 32070
rect 3329 32011 3387 32017
rect 3329 31977 3341 32011
rect 3375 32008 3387 32011
rect 3970 32008 3976 32020
rect 3375 31980 3976 32008
rect 3375 31977 3387 31980
rect 3329 31971 3387 31977
rect 3970 31968 3976 31980
rect 4028 31968 4034 32020
rect 5626 31968 5632 32020
rect 5684 32008 5690 32020
rect 5721 32011 5779 32017
rect 5721 32008 5733 32011
rect 5684 31980 5733 32008
rect 5684 31968 5690 31980
rect 5721 31977 5733 31980
rect 5767 31977 5779 32011
rect 5721 31971 5779 31977
rect 7374 31968 7380 32020
rect 7432 32008 7438 32020
rect 7837 32011 7895 32017
rect 7837 32008 7849 32011
rect 7432 31980 7849 32008
rect 7432 31968 7438 31980
rect 7837 31977 7849 31980
rect 7883 31977 7895 32011
rect 9582 32008 9588 32020
rect 9543 31980 9588 32008
rect 7837 31971 7895 31977
rect 9582 31968 9588 31980
rect 9640 31968 9646 32020
rect 10226 32008 10232 32020
rect 10187 31980 10232 32008
rect 10226 31968 10232 31980
rect 10284 31968 10290 32020
rect 12434 32008 12440 32020
rect 12395 31980 12440 32008
rect 12434 31968 12440 31980
rect 12492 31968 12498 32020
rect 12986 32008 12992 32020
rect 12947 31980 12992 32008
rect 12986 31968 12992 31980
rect 13044 31968 13050 32020
rect 15194 31968 15200 32020
rect 15252 32008 15258 32020
rect 15473 32011 15531 32017
rect 15473 32008 15485 32011
rect 15252 31980 15485 32008
rect 15252 31968 15258 31980
rect 15473 31977 15485 31980
rect 15519 31977 15531 32011
rect 15473 31971 15531 31977
rect 19981 32011 20039 32017
rect 19981 31977 19993 32011
rect 20027 32008 20039 32011
rect 20162 32008 20168 32020
rect 20027 31980 20168 32008
rect 20027 31977 20039 31980
rect 19981 31971 20039 31977
rect 20162 31968 20168 31980
rect 20220 31968 20226 32020
rect 20254 31968 20260 32020
rect 20312 32008 20318 32020
rect 20349 32011 20407 32017
rect 20349 32008 20361 32011
rect 20312 31980 20361 32008
rect 20312 31968 20318 31980
rect 20349 31977 20361 31980
rect 20395 31977 20407 32011
rect 20349 31971 20407 31977
rect 20441 32011 20499 32017
rect 20441 31977 20453 32011
rect 20487 32008 20499 32011
rect 21266 32008 21272 32020
rect 20487 31980 21272 32008
rect 20487 31977 20499 31980
rect 20441 31971 20499 31977
rect 21266 31968 21272 31980
rect 21324 31968 21330 32020
rect 26510 31968 26516 32020
rect 26568 31968 26574 32020
rect 26694 31968 26700 32020
rect 26752 32008 26758 32020
rect 27295 32011 27353 32017
rect 27295 32008 27307 32011
rect 26752 31980 27307 32008
rect 26752 31968 26758 31980
rect 27295 31977 27307 31980
rect 27341 31977 27353 32011
rect 30466 32008 30472 32020
rect 30427 31980 30472 32008
rect 27295 31971 27353 31977
rect 30466 31968 30472 31980
rect 30524 31968 30530 32020
rect 30742 31968 30748 32020
rect 30800 32008 30806 32020
rect 30837 32011 30895 32017
rect 30837 32008 30849 32011
rect 30800 31980 30849 32008
rect 30800 31968 30806 31980
rect 30837 31977 30849 31980
rect 30883 32008 30895 32011
rect 30883 31980 32168 32008
rect 30883 31977 30895 31980
rect 30837 31971 30895 31977
rect 3878 31900 3884 31952
rect 3936 31940 3942 31952
rect 6724 31943 6782 31949
rect 3936 31912 6500 31940
rect 3936 31900 3942 31912
rect 3142 31872 3148 31884
rect 3103 31844 3148 31872
rect 3142 31832 3148 31844
rect 3200 31832 3206 31884
rect 4522 31872 4528 31884
rect 4483 31844 4528 31872
rect 4522 31832 4528 31844
rect 4580 31832 4586 31884
rect 5353 31875 5411 31881
rect 5353 31841 5365 31875
rect 5399 31872 5411 31875
rect 5718 31872 5724 31884
rect 5399 31844 5724 31872
rect 5399 31841 5411 31844
rect 5353 31835 5411 31841
rect 5718 31832 5724 31844
rect 5776 31832 5782 31884
rect 6472 31881 6500 31912
rect 6724 31909 6736 31943
rect 6770 31940 6782 31943
rect 6822 31940 6828 31952
rect 6770 31912 6828 31940
rect 6770 31909 6782 31912
rect 6724 31903 6782 31909
rect 6822 31900 6828 31912
rect 6880 31900 6886 31952
rect 7282 31900 7288 31952
rect 7340 31940 7346 31952
rect 11146 31940 11152 31952
rect 7340 31912 11152 31940
rect 7340 31900 7346 31912
rect 10152 31881 10180 31912
rect 11146 31900 11152 31912
rect 11204 31940 11210 31952
rect 11204 31912 13216 31940
rect 11204 31900 11210 31912
rect 6457 31875 6515 31881
rect 6457 31841 6469 31875
rect 6503 31841 6515 31875
rect 6457 31835 6515 31841
rect 9677 31875 9735 31881
rect 9677 31841 9689 31875
rect 9723 31841 9735 31875
rect 9677 31835 9735 31841
rect 10137 31875 10195 31881
rect 10137 31841 10149 31875
rect 10183 31841 10195 31875
rect 10137 31835 10195 31841
rect 10321 31875 10379 31881
rect 10321 31841 10333 31875
rect 10367 31872 10379 31875
rect 10410 31872 10416 31884
rect 10367 31844 10416 31872
rect 10367 31841 10379 31844
rect 10321 31835 10379 31841
rect 2961 31807 3019 31813
rect 2961 31773 2973 31807
rect 3007 31804 3019 31807
rect 4338 31804 4344 31816
rect 3007 31776 4344 31804
rect 3007 31773 3019 31776
rect 2961 31767 3019 31773
rect 4338 31764 4344 31776
rect 4396 31764 4402 31816
rect 4709 31807 4767 31813
rect 4709 31773 4721 31807
rect 4755 31804 4767 31807
rect 5261 31807 5319 31813
rect 5261 31804 5273 31807
rect 4755 31776 5273 31804
rect 4755 31773 4767 31776
rect 4709 31767 4767 31773
rect 5261 31773 5273 31776
rect 5307 31773 5319 31807
rect 5442 31804 5448 31816
rect 5403 31776 5448 31804
rect 5261 31767 5319 31773
rect 5442 31764 5448 31776
rect 5500 31764 5506 31816
rect 5537 31807 5595 31813
rect 5537 31773 5549 31807
rect 5583 31773 5595 31807
rect 9692 31804 9720 31835
rect 10410 31832 10416 31844
rect 10468 31832 10474 31884
rect 12360 31881 12388 31912
rect 13188 31881 13216 31912
rect 14366 31900 14372 31952
rect 14424 31940 14430 31952
rect 15013 31943 15071 31949
rect 15013 31940 15025 31943
rect 14424 31912 15025 31940
rect 14424 31900 14430 31912
rect 15013 31909 15025 31912
rect 15059 31909 15071 31943
rect 15013 31903 15071 31909
rect 17402 31900 17408 31952
rect 17460 31900 17466 31952
rect 21910 31900 21916 31952
rect 21968 31940 21974 31952
rect 21968 31912 22126 31940
rect 26528 31926 26556 31968
rect 29089 31943 29147 31949
rect 21968 31900 21974 31912
rect 29089 31909 29101 31943
rect 29135 31940 29147 31943
rect 29270 31940 29276 31952
rect 29135 31912 29276 31940
rect 29135 31909 29147 31912
rect 29089 31903 29147 31909
rect 29270 31900 29276 31912
rect 29328 31940 29334 31952
rect 30006 31940 30012 31952
rect 29328 31912 30012 31940
rect 29328 31900 29334 31912
rect 30006 31900 30012 31912
rect 30064 31900 30070 31952
rect 32140 31949 32168 31980
rect 32125 31943 32183 31949
rect 32125 31909 32137 31943
rect 32171 31909 32183 31943
rect 32125 31903 32183 31909
rect 12345 31875 12403 31881
rect 12345 31841 12357 31875
rect 12391 31841 12403 31875
rect 12345 31835 12403 31841
rect 12989 31875 13047 31881
rect 12989 31841 13001 31875
rect 13035 31841 13047 31875
rect 12989 31835 13047 31841
rect 13173 31875 13231 31881
rect 13173 31841 13185 31875
rect 13219 31841 13231 31875
rect 15102 31872 15108 31884
rect 15063 31844 15108 31872
rect 13173 31835 13231 31841
rect 9858 31804 9864 31816
rect 9692 31776 9864 31804
rect 5537 31767 5595 31773
rect 5552 31736 5580 31767
rect 9858 31764 9864 31776
rect 9916 31804 9922 31816
rect 13004 31804 13032 31835
rect 15102 31832 15108 31844
rect 15160 31832 15166 31884
rect 16209 31875 16267 31881
rect 16209 31841 16221 31875
rect 16255 31872 16267 31875
rect 16298 31872 16304 31884
rect 16255 31844 16304 31872
rect 16255 31841 16267 31844
rect 16209 31835 16267 31841
rect 16298 31832 16304 31844
rect 16356 31832 16362 31884
rect 23014 31832 23020 31884
rect 23072 31872 23078 31884
rect 23109 31875 23167 31881
rect 23109 31872 23121 31875
rect 23072 31844 23121 31872
rect 23072 31832 23078 31844
rect 23109 31841 23121 31844
rect 23155 31841 23167 31875
rect 25866 31872 25872 31884
rect 25827 31844 25872 31872
rect 23109 31835 23167 31841
rect 25866 31832 25872 31844
rect 25924 31832 25930 31884
rect 28997 31875 29055 31881
rect 28997 31841 29009 31875
rect 29043 31872 29055 31875
rect 29546 31872 29552 31884
rect 29043 31844 29552 31872
rect 29043 31841 29055 31844
rect 28997 31835 29055 31841
rect 29546 31832 29552 31844
rect 29604 31832 29610 31884
rect 29840 31844 31156 31872
rect 9916 31776 13032 31804
rect 14829 31807 14887 31813
rect 9916 31764 9922 31776
rect 14829 31773 14841 31807
rect 14875 31773 14887 31807
rect 14829 31767 14887 31773
rect 5718 31736 5724 31748
rect 5552 31708 5724 31736
rect 5718 31696 5724 31708
rect 5776 31696 5782 31748
rect 9674 31696 9680 31748
rect 9732 31736 9738 31748
rect 10042 31736 10048 31748
rect 9732 31708 10048 31736
rect 9732 31696 9738 31708
rect 10042 31696 10048 31708
rect 10100 31696 10106 31748
rect 12802 31736 12808 31748
rect 12406 31708 12808 31736
rect 7190 31628 7196 31680
rect 7248 31668 7254 31680
rect 12406 31668 12434 31708
rect 12802 31696 12808 31708
rect 12860 31736 12866 31748
rect 13170 31736 13176 31748
rect 12860 31708 13176 31736
rect 12860 31696 12866 31708
rect 13170 31696 13176 31708
rect 13228 31696 13234 31748
rect 7248 31640 12434 31668
rect 7248 31628 7254 31640
rect 12526 31628 12532 31680
rect 12584 31668 12590 31680
rect 14844 31668 14872 31767
rect 16574 31764 16580 31816
rect 16632 31804 16638 31816
rect 20625 31807 20683 31813
rect 16632 31776 16677 31804
rect 16632 31764 16638 31776
rect 20625 31773 20637 31807
rect 20671 31773 20683 31807
rect 20625 31767 20683 31773
rect 21683 31807 21741 31813
rect 21683 31773 21695 31807
rect 21729 31804 21741 31807
rect 22094 31804 22100 31816
rect 21729 31776 22100 31804
rect 21729 31773 21741 31776
rect 21683 31767 21741 31773
rect 20640 31736 20668 31767
rect 22094 31764 22100 31776
rect 22152 31764 22158 31816
rect 23477 31807 23535 31813
rect 23477 31773 23489 31807
rect 23523 31804 23535 31807
rect 23566 31804 23572 31816
rect 23523 31776 23572 31804
rect 23523 31773 23535 31776
rect 23477 31767 23535 31773
rect 23566 31764 23572 31776
rect 23624 31804 23630 31816
rect 25501 31807 25559 31813
rect 25501 31804 25513 31807
rect 23624 31776 25513 31804
rect 23624 31764 23630 31776
rect 25501 31773 25513 31776
rect 25547 31773 25559 31807
rect 25501 31767 25559 31773
rect 29273 31807 29331 31813
rect 29273 31773 29285 31807
rect 29319 31804 29331 31807
rect 29454 31804 29460 31816
rect 29319 31776 29460 31804
rect 29319 31773 29331 31776
rect 29273 31767 29331 31773
rect 29454 31764 29460 31776
rect 29512 31804 29518 31816
rect 29840 31804 29868 31844
rect 29512 31776 29868 31804
rect 29512 31764 29518 31776
rect 29914 31764 29920 31816
rect 29972 31804 29978 31816
rect 31128 31813 31156 31844
rect 30929 31807 30987 31813
rect 29972 31776 30880 31804
rect 29972 31764 29978 31776
rect 20714 31736 20720 31748
rect 20640 31708 20720 31736
rect 20714 31696 20720 31708
rect 20772 31696 20778 31748
rect 29362 31696 29368 31748
rect 29420 31736 29426 31748
rect 30650 31736 30656 31748
rect 29420 31708 30656 31736
rect 29420 31696 29426 31708
rect 30650 31696 30656 31708
rect 30708 31696 30714 31748
rect 12584 31640 14872 31668
rect 12584 31628 12590 31640
rect 17954 31628 17960 31680
rect 18012 31677 18018 31680
rect 18012 31671 18061 31677
rect 18012 31637 18015 31671
rect 18049 31637 18061 31671
rect 18012 31631 18061 31637
rect 18012 31628 18018 31631
rect 28074 31628 28080 31680
rect 28132 31668 28138 31680
rect 28629 31671 28687 31677
rect 28629 31668 28641 31671
rect 28132 31640 28641 31668
rect 28132 31628 28138 31640
rect 28629 31637 28641 31640
rect 28675 31637 28687 31671
rect 30852 31668 30880 31776
rect 30929 31773 30941 31807
rect 30975 31773 30987 31807
rect 30929 31767 30987 31773
rect 31113 31807 31171 31813
rect 31113 31773 31125 31807
rect 31159 31804 31171 31807
rect 31202 31804 31208 31816
rect 31159 31776 31208 31804
rect 31159 31773 31171 31776
rect 31113 31767 31171 31773
rect 30944 31736 30972 31767
rect 31202 31764 31208 31776
rect 31260 31764 31266 31816
rect 31662 31764 31668 31816
rect 31720 31764 31726 31816
rect 31680 31736 31708 31764
rect 31757 31739 31815 31745
rect 31757 31736 31769 31739
rect 30944 31708 31769 31736
rect 31757 31705 31769 31708
rect 31803 31705 31815 31739
rect 31757 31699 31815 31705
rect 31665 31671 31723 31677
rect 31665 31668 31677 31671
rect 30852 31640 31677 31668
rect 28629 31631 28687 31637
rect 31665 31637 31677 31640
rect 31711 31637 31723 31671
rect 31665 31631 31723 31637
rect 1104 31578 34316 31600
rect 1104 31526 6517 31578
rect 6569 31526 6581 31578
rect 6633 31526 6645 31578
rect 6697 31526 6709 31578
rect 6761 31526 17588 31578
rect 17640 31526 17652 31578
rect 17704 31526 17716 31578
rect 17768 31526 17780 31578
rect 17832 31526 28658 31578
rect 28710 31526 28722 31578
rect 28774 31526 28786 31578
rect 28838 31526 28850 31578
rect 28902 31526 34316 31578
rect 1104 31504 34316 31526
rect 13909 31467 13967 31473
rect 4172 31436 10364 31464
rect 3142 31288 3148 31340
rect 3200 31328 3206 31340
rect 3694 31328 3700 31340
rect 3200 31300 3700 31328
rect 3200 31288 3206 31300
rect 3694 31288 3700 31300
rect 3752 31328 3758 31340
rect 4065 31331 4123 31337
rect 4065 31328 4077 31331
rect 3752 31300 4077 31328
rect 3752 31288 3758 31300
rect 4065 31297 4077 31300
rect 4111 31297 4123 31331
rect 4065 31291 4123 31297
rect 3973 31263 4031 31269
rect 3973 31229 3985 31263
rect 4019 31260 4031 31263
rect 4172 31260 4200 31436
rect 4338 31356 4344 31408
rect 4396 31396 4402 31408
rect 4396 31368 6868 31396
rect 4396 31356 4402 31368
rect 4249 31331 4307 31337
rect 4249 31297 4261 31331
rect 4295 31328 4307 31331
rect 4982 31328 4988 31340
rect 4295 31300 4988 31328
rect 4295 31297 4307 31300
rect 4249 31291 4307 31297
rect 4982 31288 4988 31300
rect 5040 31328 5046 31340
rect 5350 31328 5356 31340
rect 5040 31300 5356 31328
rect 5040 31288 5046 31300
rect 5350 31288 5356 31300
rect 5408 31288 5414 31340
rect 4019 31232 4200 31260
rect 4019 31229 4031 31232
rect 3973 31223 4031 31229
rect 5534 31220 5540 31272
rect 5592 31260 5598 31272
rect 6840 31269 6868 31368
rect 5629 31263 5687 31269
rect 5629 31260 5641 31263
rect 5592 31232 5641 31260
rect 5592 31220 5598 31232
rect 5629 31229 5641 31232
rect 5675 31229 5687 31263
rect 5629 31223 5687 31229
rect 5905 31263 5963 31269
rect 5905 31229 5917 31263
rect 5951 31229 5963 31263
rect 5905 31223 5963 31229
rect 6825 31263 6883 31269
rect 6825 31229 6837 31263
rect 6871 31229 6883 31263
rect 6825 31223 6883 31229
rect 7009 31263 7067 31269
rect 7009 31229 7021 31263
rect 7055 31260 7067 31263
rect 7374 31260 7380 31272
rect 7055 31232 7380 31260
rect 7055 31229 7067 31232
rect 7009 31223 7067 31229
rect 5920 31192 5948 31223
rect 7024 31192 7052 31223
rect 7374 31220 7380 31232
rect 7432 31220 7438 31272
rect 9493 31263 9551 31269
rect 9493 31229 9505 31263
rect 9539 31260 9551 31263
rect 9950 31260 9956 31272
rect 9539 31232 9956 31260
rect 9539 31229 9551 31232
rect 9493 31223 9551 31229
rect 9950 31220 9956 31232
rect 10008 31220 10014 31272
rect 10336 31269 10364 31436
rect 13909 31433 13921 31467
rect 13955 31464 13967 31467
rect 15102 31464 15108 31476
rect 13955 31436 15108 31464
rect 13955 31433 13967 31436
rect 13909 31427 13967 31433
rect 15102 31424 15108 31436
rect 15160 31424 15166 31476
rect 16574 31424 16580 31476
rect 16632 31464 16638 31476
rect 17497 31467 17555 31473
rect 17497 31464 17509 31467
rect 16632 31436 17509 31464
rect 16632 31424 16638 31436
rect 17497 31433 17509 31436
rect 17543 31433 17555 31467
rect 17497 31427 17555 31433
rect 20714 31424 20720 31476
rect 20772 31464 20778 31476
rect 22649 31467 22707 31473
rect 22649 31464 22661 31467
rect 20772 31436 22661 31464
rect 20772 31424 20778 31436
rect 22649 31433 22661 31436
rect 22695 31433 22707 31467
rect 22649 31427 22707 31433
rect 18969 31399 19027 31405
rect 18969 31396 18981 31399
rect 17788 31368 18981 31396
rect 12526 31328 12532 31340
rect 12487 31300 12532 31328
rect 12526 31288 12532 31300
rect 12584 31288 12590 31340
rect 10137 31263 10195 31269
rect 10137 31229 10149 31263
rect 10183 31229 10195 31263
rect 10137 31223 10195 31229
rect 10321 31263 10379 31269
rect 10321 31229 10333 31263
rect 10367 31260 10379 31263
rect 11606 31260 11612 31272
rect 10367 31232 11612 31260
rect 10367 31229 10379 31232
rect 10321 31223 10379 31229
rect 5920 31164 7052 31192
rect 9248 31195 9306 31201
rect 9248 31161 9260 31195
rect 9294 31192 9306 31195
rect 9766 31192 9772 31204
rect 9294 31164 9772 31192
rect 9294 31161 9306 31164
rect 9248 31155 9306 31161
rect 9766 31152 9772 31164
rect 9824 31152 9830 31204
rect 9858 31152 9864 31204
rect 9916 31192 9922 31204
rect 10152 31192 10180 31223
rect 11606 31220 11612 31232
rect 11664 31260 11670 31272
rect 12621 31263 12679 31269
rect 12621 31260 12633 31263
rect 11664 31232 12633 31260
rect 11664 31220 11670 31232
rect 12621 31229 12633 31232
rect 12667 31229 12679 31263
rect 12621 31223 12679 31229
rect 13354 31220 13360 31272
rect 13412 31260 13418 31272
rect 13725 31263 13783 31269
rect 13725 31260 13737 31263
rect 13412 31232 13737 31260
rect 13412 31220 13418 31232
rect 13725 31229 13737 31232
rect 13771 31229 13783 31263
rect 13906 31260 13912 31272
rect 13867 31232 13912 31260
rect 13725 31223 13783 31229
rect 13906 31220 13912 31232
rect 13964 31220 13970 31272
rect 15749 31263 15807 31269
rect 15749 31229 15761 31263
rect 15795 31260 15807 31263
rect 16114 31260 16120 31272
rect 15795 31232 16120 31260
rect 15795 31229 15807 31232
rect 15749 31223 15807 31229
rect 16114 31220 16120 31232
rect 16172 31220 16178 31272
rect 9916 31164 10180 31192
rect 9916 31152 9922 31164
rect 15286 31152 15292 31204
rect 15344 31192 15350 31204
rect 15482 31195 15540 31201
rect 15482 31192 15494 31195
rect 15344 31164 15494 31192
rect 15344 31152 15350 31164
rect 15482 31161 15494 31164
rect 15528 31161 15540 31195
rect 17788 31192 17816 31368
rect 18969 31365 18981 31368
rect 19015 31365 19027 31399
rect 18969 31359 19027 31365
rect 18138 31328 18144 31340
rect 18099 31300 18144 31328
rect 18138 31288 18144 31300
rect 18196 31288 18202 31340
rect 18598 31288 18604 31340
rect 18656 31328 18662 31340
rect 18840 31331 18898 31337
rect 18840 31328 18852 31331
rect 18656 31300 18852 31328
rect 18656 31288 18662 31300
rect 18840 31297 18852 31300
rect 18886 31297 18898 31331
rect 18840 31291 18898 31297
rect 19061 31331 19119 31337
rect 19061 31297 19073 31331
rect 19107 31297 19119 31331
rect 23566 31328 23572 31340
rect 23527 31300 23572 31328
rect 19061 31291 19119 31297
rect 17954 31260 17960 31272
rect 17867 31232 17960 31260
rect 17954 31220 17960 31232
rect 18012 31260 18018 31272
rect 19076 31260 19104 31291
rect 23566 31288 23572 31300
rect 23624 31288 23630 31340
rect 24302 31288 24308 31340
rect 24360 31328 24366 31340
rect 28074 31328 28080 31340
rect 24360 31300 24992 31328
rect 28035 31300 28080 31328
rect 24360 31288 24366 31300
rect 22830 31260 22836 31272
rect 18012 31232 19104 31260
rect 22791 31232 22836 31260
rect 18012 31220 18018 31232
rect 22830 31220 22836 31232
rect 22888 31220 22894 31272
rect 23934 31260 23940 31272
rect 23895 31232 23940 31260
rect 23934 31220 23940 31232
rect 23992 31220 23998 31272
rect 17865 31195 17923 31201
rect 17865 31192 17877 31195
rect 17788 31164 17877 31192
rect 15482 31155 15540 31161
rect 17865 31161 17877 31164
rect 17911 31161 17923 31195
rect 17865 31155 17923 31161
rect 18693 31195 18751 31201
rect 18693 31161 18705 31195
rect 18739 31192 18751 31195
rect 19610 31192 19616 31204
rect 18739 31164 19616 31192
rect 18739 31161 18751 31164
rect 18693 31155 18751 31161
rect 3142 31084 3148 31136
rect 3200 31124 3206 31136
rect 3605 31127 3663 31133
rect 3605 31124 3617 31127
rect 3200 31096 3617 31124
rect 3200 31084 3206 31096
rect 3605 31093 3617 31096
rect 3651 31093 3663 31127
rect 3605 31087 3663 31093
rect 5813 31127 5871 31133
rect 5813 31093 5825 31127
rect 5859 31124 5871 31127
rect 5902 31124 5908 31136
rect 5859 31096 5908 31124
rect 5859 31093 5871 31096
rect 5813 31087 5871 31093
rect 5902 31084 5908 31096
rect 5960 31084 5966 31136
rect 7098 31084 7104 31136
rect 7156 31124 7162 31136
rect 7193 31127 7251 31133
rect 7193 31124 7205 31127
rect 7156 31096 7205 31124
rect 7156 31084 7162 31096
rect 7193 31093 7205 31096
rect 7239 31093 7251 31127
rect 7193 31087 7251 31093
rect 8113 31127 8171 31133
rect 8113 31093 8125 31127
rect 8159 31124 8171 31127
rect 8202 31124 8208 31136
rect 8159 31096 8208 31124
rect 8159 31093 8171 31096
rect 8113 31087 8171 31093
rect 8202 31084 8208 31096
rect 8260 31084 8266 31136
rect 10134 31124 10140 31136
rect 10095 31096 10140 31124
rect 10134 31084 10140 31096
rect 10192 31084 10198 31136
rect 12434 31084 12440 31136
rect 12492 31124 12498 31136
rect 12713 31127 12771 31133
rect 12713 31124 12725 31127
rect 12492 31096 12725 31124
rect 12492 31084 12498 31096
rect 12713 31093 12725 31096
rect 12759 31093 12771 31127
rect 13078 31124 13084 31136
rect 13039 31096 13084 31124
rect 12713 31087 12771 31093
rect 13078 31084 13084 31096
rect 13136 31084 13142 31136
rect 14366 31124 14372 31136
rect 14327 31096 14372 31124
rect 14366 31084 14372 31096
rect 14424 31084 14430 31136
rect 17880 31124 17908 31155
rect 19610 31152 19616 31164
rect 19668 31152 19674 31204
rect 24964 31192 24992 31300
rect 28074 31288 28080 31300
rect 28132 31288 28138 31340
rect 31294 31288 31300 31340
rect 31352 31328 31358 31340
rect 31389 31331 31447 31337
rect 31389 31328 31401 31331
rect 31352 31300 31401 31328
rect 31352 31288 31358 31300
rect 31389 31297 31401 31300
rect 31435 31297 31447 31331
rect 31389 31291 31447 31297
rect 27614 31220 27620 31272
rect 27672 31260 27678 31272
rect 27798 31260 27804 31272
rect 27672 31232 27804 31260
rect 27672 31220 27678 31232
rect 27798 31220 27804 31232
rect 27856 31220 27862 31272
rect 31205 31263 31263 31269
rect 31205 31229 31217 31263
rect 31251 31260 31263 31263
rect 31662 31260 31668 31272
rect 31251 31232 31668 31260
rect 31251 31229 31263 31232
rect 31205 31223 31263 31229
rect 31662 31220 31668 31232
rect 31720 31220 31726 31272
rect 26510 31192 26516 31204
rect 24964 31178 26516 31192
rect 24978 31164 26516 31178
rect 26510 31152 26516 31164
rect 26568 31152 26574 31204
rect 29362 31192 29368 31204
rect 29302 31164 29368 31192
rect 29362 31152 29368 31164
rect 29420 31152 29426 31204
rect 17954 31124 17960 31136
rect 17880 31096 17960 31124
rect 17954 31084 17960 31096
rect 18012 31084 18018 31136
rect 19058 31084 19064 31136
rect 19116 31124 19122 31136
rect 19337 31127 19395 31133
rect 19337 31124 19349 31127
rect 19116 31096 19349 31124
rect 19116 31084 19122 31096
rect 19337 31093 19349 31096
rect 19383 31093 19395 31127
rect 19337 31087 19395 31093
rect 25314 31084 25320 31136
rect 25372 31133 25378 31136
rect 25372 31127 25421 31133
rect 25372 31093 25375 31127
rect 25409 31093 25421 31127
rect 29546 31124 29552 31136
rect 29507 31096 29552 31124
rect 25372 31087 25421 31093
rect 25372 31084 25378 31087
rect 29546 31084 29552 31096
rect 29604 31084 29610 31136
rect 30837 31127 30895 31133
rect 30837 31093 30849 31127
rect 30883 31124 30895 31127
rect 31018 31124 31024 31136
rect 30883 31096 31024 31124
rect 30883 31093 30895 31096
rect 30837 31087 30895 31093
rect 31018 31084 31024 31096
rect 31076 31084 31082 31136
rect 31294 31124 31300 31136
rect 31255 31096 31300 31124
rect 31294 31084 31300 31096
rect 31352 31084 31358 31136
rect 1104 31034 34316 31056
rect 1104 30982 12052 31034
rect 12104 30982 12116 31034
rect 12168 30982 12180 31034
rect 12232 30982 12244 31034
rect 12296 30982 23123 31034
rect 23175 30982 23187 31034
rect 23239 30982 23251 31034
rect 23303 30982 23315 31034
rect 23367 30982 34316 31034
rect 1104 30960 34316 30982
rect 6641 30923 6699 30929
rect 6641 30889 6653 30923
rect 6687 30920 6699 30923
rect 6822 30920 6828 30932
rect 6687 30892 6828 30920
rect 6687 30889 6699 30892
rect 6641 30883 6699 30889
rect 6822 30880 6828 30892
rect 6880 30880 6886 30932
rect 11606 30920 11612 30932
rect 11567 30892 11612 30920
rect 11606 30880 11612 30892
rect 11664 30880 11670 30932
rect 12434 30880 12440 30932
rect 12492 30920 12498 30932
rect 12492 30892 12537 30920
rect 12492 30880 12498 30892
rect 13906 30880 13912 30932
rect 13964 30920 13970 30932
rect 14829 30923 14887 30929
rect 14829 30920 14841 30923
rect 13964 30892 14841 30920
rect 13964 30880 13970 30892
rect 14829 30889 14841 30892
rect 14875 30920 14887 30923
rect 14918 30920 14924 30932
rect 14875 30892 14924 30920
rect 14875 30889 14887 30892
rect 14829 30883 14887 30889
rect 14918 30880 14924 30892
rect 14976 30880 14982 30932
rect 17954 30929 17960 30932
rect 17911 30923 17960 30929
rect 17911 30889 17923 30923
rect 17957 30889 17960 30923
rect 17911 30883 17960 30889
rect 17954 30880 17960 30883
rect 18012 30880 18018 30932
rect 23017 30923 23075 30929
rect 23017 30889 23029 30923
rect 23063 30920 23075 30923
rect 23474 30920 23480 30932
rect 23063 30892 23480 30920
rect 23063 30889 23075 30892
rect 23017 30883 23075 30889
rect 23474 30880 23480 30892
rect 23532 30880 23538 30932
rect 23569 30923 23627 30929
rect 23569 30889 23581 30923
rect 23615 30920 23627 30923
rect 23934 30920 23940 30932
rect 23615 30892 23940 30920
rect 23615 30889 23627 30892
rect 23569 30883 23627 30889
rect 23934 30880 23940 30892
rect 23992 30880 23998 30932
rect 24029 30923 24087 30929
rect 24029 30889 24041 30923
rect 24075 30920 24087 30923
rect 25314 30920 25320 30932
rect 24075 30892 25320 30920
rect 24075 30889 24087 30892
rect 24029 30883 24087 30889
rect 25314 30880 25320 30892
rect 25372 30880 25378 30932
rect 30650 30880 30656 30932
rect 30708 30920 30714 30932
rect 30708 30892 31524 30920
rect 30708 30880 30714 30892
rect 5442 30812 5448 30864
rect 5500 30852 5506 30864
rect 11624 30852 11652 30880
rect 12805 30855 12863 30861
rect 12805 30852 12817 30855
rect 5500 30824 6960 30852
rect 11624 30824 12817 30852
rect 5500 30812 5506 30824
rect 3142 30784 3148 30796
rect 3103 30756 3148 30784
rect 3142 30744 3148 30756
rect 3200 30744 3206 30796
rect 4798 30744 4804 30796
rect 4856 30784 4862 30796
rect 5261 30787 5319 30793
rect 5261 30784 5273 30787
rect 4856 30756 5273 30784
rect 4856 30744 4862 30756
rect 5261 30753 5273 30756
rect 5307 30753 5319 30787
rect 5626 30784 5632 30796
rect 5587 30756 5632 30784
rect 5261 30747 5319 30753
rect 5626 30744 5632 30756
rect 5684 30744 5690 30796
rect 5902 30784 5908 30796
rect 5863 30756 5908 30784
rect 5902 30744 5908 30756
rect 5960 30744 5966 30796
rect 6932 30793 6960 30824
rect 12805 30821 12817 30824
rect 12851 30821 12863 30855
rect 12805 30815 12863 30821
rect 17402 30812 17408 30864
rect 17460 30812 17466 30864
rect 23492 30852 23520 30880
rect 31496 30864 31524 30892
rect 31662 30880 31668 30932
rect 31720 30920 31726 30932
rect 32493 30923 32551 30929
rect 32493 30920 32505 30923
rect 31720 30892 32505 30920
rect 31720 30880 31726 30892
rect 32493 30889 32505 30892
rect 32539 30889 32551 30923
rect 32493 30883 32551 30889
rect 23492 30824 24072 30852
rect 6917 30787 6975 30793
rect 6917 30753 6929 30787
rect 6963 30753 6975 30787
rect 7098 30784 7104 30796
rect 7059 30756 7104 30784
rect 6917 30747 6975 30753
rect 7098 30744 7104 30756
rect 7156 30744 7162 30796
rect 10042 30744 10048 30796
rect 10100 30784 10106 30796
rect 10485 30787 10543 30793
rect 10485 30784 10497 30787
rect 10100 30756 10497 30784
rect 10100 30744 10106 30756
rect 10485 30753 10497 30756
rect 10531 30753 10543 30787
rect 10485 30747 10543 30753
rect 12618 30744 12624 30796
rect 12676 30784 12682 30796
rect 12897 30787 12955 30793
rect 12897 30784 12909 30787
rect 12676 30756 12909 30784
rect 12676 30744 12682 30756
rect 12897 30753 12909 30756
rect 12943 30784 12955 30787
rect 13630 30784 13636 30796
rect 12943 30756 13636 30784
rect 12943 30753 12955 30756
rect 12897 30747 12955 30753
rect 13630 30744 13636 30756
rect 13688 30744 13694 30796
rect 14366 30744 14372 30796
rect 14424 30784 14430 30796
rect 14737 30787 14795 30793
rect 14737 30784 14749 30787
rect 14424 30756 14749 30784
rect 14424 30744 14430 30756
rect 14737 30753 14749 30756
rect 14783 30753 14795 30787
rect 20530 30784 20536 30796
rect 20491 30756 20536 30784
rect 14737 30747 14795 30753
rect 20530 30744 20536 30756
rect 20588 30744 20594 30796
rect 22830 30784 22836 30796
rect 22743 30756 22836 30784
rect 22830 30744 22836 30756
rect 22888 30784 22894 30796
rect 23934 30784 23940 30796
rect 22888 30756 23152 30784
rect 23895 30756 23940 30784
rect 22888 30744 22894 30756
rect 2958 30716 2964 30728
rect 2871 30688 2964 30716
rect 2958 30676 2964 30688
rect 3016 30676 3022 30728
rect 3050 30676 3056 30728
rect 3108 30716 3114 30728
rect 3234 30716 3240 30728
rect 3108 30688 3153 30716
rect 3195 30688 3240 30716
rect 3108 30676 3114 30688
rect 3234 30676 3240 30688
rect 3292 30676 3298 30728
rect 4982 30716 4988 30728
rect 4943 30688 4988 30716
rect 4982 30676 4988 30688
rect 5040 30676 5046 30728
rect 6825 30719 6883 30725
rect 6825 30685 6837 30719
rect 6871 30685 6883 30719
rect 7006 30716 7012 30728
rect 6967 30688 7012 30716
rect 6825 30679 6883 30685
rect 2774 30540 2780 30592
rect 2832 30580 2838 30592
rect 2976 30580 3004 30676
rect 4062 30608 4068 30660
rect 4120 30648 4126 30660
rect 5718 30648 5724 30660
rect 4120 30620 5724 30648
rect 4120 30608 4126 30620
rect 5718 30608 5724 30620
rect 5776 30648 5782 30660
rect 6840 30648 6868 30679
rect 7006 30676 7012 30688
rect 7064 30676 7070 30728
rect 9950 30676 9956 30728
rect 10008 30716 10014 30728
rect 10229 30719 10287 30725
rect 10229 30716 10241 30719
rect 10008 30688 10241 30716
rect 10008 30676 10014 30688
rect 10229 30685 10241 30688
rect 10275 30685 10287 30719
rect 10229 30679 10287 30685
rect 13081 30719 13139 30725
rect 13081 30685 13093 30719
rect 13127 30716 13139 30719
rect 13354 30716 13360 30728
rect 13127 30688 13360 30716
rect 13127 30685 13139 30688
rect 13081 30679 13139 30685
rect 5776 30620 6868 30648
rect 5776 30608 5782 30620
rect 4080 30580 4108 30608
rect 2832 30552 2877 30580
rect 2976 30552 4108 30580
rect 10244 30580 10272 30679
rect 13354 30676 13360 30688
rect 13412 30676 13418 30728
rect 16114 30716 16120 30728
rect 16075 30688 16120 30716
rect 16114 30676 16120 30688
rect 16172 30676 16178 30728
rect 16485 30719 16543 30725
rect 16485 30685 16497 30719
rect 16531 30716 16543 30719
rect 17402 30716 17408 30728
rect 16531 30688 17408 30716
rect 16531 30685 16543 30688
rect 16485 30679 16543 30685
rect 17402 30676 17408 30688
rect 17460 30676 17466 30728
rect 19610 30676 19616 30728
rect 19668 30716 19674 30728
rect 20625 30719 20683 30725
rect 20625 30716 20637 30719
rect 19668 30688 20637 30716
rect 19668 30676 19674 30688
rect 20625 30685 20637 30688
rect 20671 30685 20683 30719
rect 20625 30679 20683 30685
rect 20717 30719 20775 30725
rect 20717 30685 20729 30719
rect 20763 30685 20775 30719
rect 20717 30679 20775 30685
rect 20346 30608 20352 30660
rect 20404 30648 20410 30660
rect 20732 30648 20760 30679
rect 20404 30620 20760 30648
rect 23124 30648 23152 30756
rect 23934 30744 23940 30756
rect 23992 30744 23998 30796
rect 24044 30784 24072 30824
rect 26510 30812 26516 30864
rect 26568 30812 26574 30864
rect 31018 30852 31024 30864
rect 30979 30824 31024 30852
rect 31018 30812 31024 30824
rect 31076 30812 31082 30864
rect 31478 30812 31484 30864
rect 31536 30812 31542 30864
rect 24044 30756 24164 30784
rect 24136 30725 24164 30756
rect 27614 30744 27620 30796
rect 27672 30784 27678 30796
rect 27709 30787 27767 30793
rect 27709 30784 27721 30787
rect 27672 30756 27721 30784
rect 27672 30744 27678 30756
rect 27709 30753 27721 30756
rect 27755 30784 27767 30787
rect 30745 30787 30803 30793
rect 30745 30784 30757 30787
rect 27755 30756 30757 30784
rect 27755 30753 27767 30756
rect 27709 30747 27767 30753
rect 30745 30753 30757 30756
rect 30791 30753 30803 30787
rect 30745 30747 30803 30753
rect 24121 30719 24179 30725
rect 24121 30685 24133 30719
rect 24167 30685 24179 30719
rect 24121 30679 24179 30685
rect 25915 30719 25973 30725
rect 25915 30685 25927 30719
rect 25961 30716 25973 30719
rect 26234 30716 26240 30728
rect 25961 30688 26240 30716
rect 25961 30685 25973 30688
rect 25915 30679 25973 30685
rect 26234 30676 26240 30688
rect 26292 30676 26298 30728
rect 27338 30716 27344 30728
rect 27299 30688 27344 30716
rect 27338 30676 27344 30688
rect 27396 30676 27402 30728
rect 24854 30648 24860 30660
rect 23124 30620 24860 30648
rect 20404 30608 20410 30620
rect 24854 30608 24860 30620
rect 24912 30608 24918 30660
rect 10870 30580 10876 30592
rect 10244 30552 10876 30580
rect 2832 30540 2838 30552
rect 10870 30540 10876 30552
rect 10928 30540 10934 30592
rect 20165 30583 20223 30589
rect 20165 30549 20177 30583
rect 20211 30580 20223 30583
rect 21082 30580 21088 30592
rect 20211 30552 21088 30580
rect 20211 30549 20223 30552
rect 20165 30543 20223 30549
rect 21082 30540 21088 30552
rect 21140 30540 21146 30592
rect 1104 30490 34316 30512
rect 1104 30438 6517 30490
rect 6569 30438 6581 30490
rect 6633 30438 6645 30490
rect 6697 30438 6709 30490
rect 6761 30438 17588 30490
rect 17640 30438 17652 30490
rect 17704 30438 17716 30490
rect 17768 30438 17780 30490
rect 17832 30438 28658 30490
rect 28710 30438 28722 30490
rect 28774 30438 28786 30490
rect 28838 30438 28850 30490
rect 28902 30438 34316 30490
rect 1104 30416 34316 30438
rect 4798 30336 4804 30388
rect 4856 30376 4862 30388
rect 10042 30376 10048 30388
rect 4856 30348 4901 30376
rect 10003 30348 10048 30376
rect 4856 30336 4862 30348
rect 10042 30336 10048 30348
rect 10100 30336 10106 30388
rect 23566 30376 23572 30388
rect 13648 30348 13860 30376
rect 6825 30311 6883 30317
rect 6825 30277 6837 30311
rect 6871 30308 6883 30311
rect 7006 30308 7012 30320
rect 6871 30280 7012 30308
rect 6871 30277 6883 30280
rect 6825 30271 6883 30277
rect 7006 30268 7012 30280
rect 7064 30268 7070 30320
rect 13173 30311 13231 30317
rect 13173 30277 13185 30311
rect 13219 30308 13231 30311
rect 13648 30308 13676 30348
rect 13219 30280 13676 30308
rect 13725 30311 13783 30317
rect 13219 30277 13231 30280
rect 13173 30271 13231 30277
rect 13725 30277 13737 30311
rect 13771 30277 13783 30311
rect 13832 30308 13860 30348
rect 22664 30348 23572 30376
rect 15105 30311 15163 30317
rect 13832 30280 14412 30308
rect 13725 30271 13783 30277
rect 7466 30240 7472 30252
rect 7427 30212 7472 30240
rect 7466 30200 7472 30212
rect 7524 30200 7530 30252
rect 10612 30212 13032 30240
rect 10612 30184 10640 30212
rect 13004 30184 13032 30212
rect 1394 30172 1400 30184
rect 1355 30144 1400 30172
rect 1394 30132 1400 30144
rect 1452 30132 1458 30184
rect 1664 30175 1722 30181
rect 1664 30141 1676 30175
rect 1710 30172 1722 30175
rect 2774 30172 2780 30184
rect 1710 30144 2780 30172
rect 1710 30141 1722 30144
rect 1664 30135 1722 30141
rect 2774 30132 2780 30144
rect 2832 30132 2838 30184
rect 3694 30172 3700 30184
rect 3655 30144 3700 30172
rect 3694 30132 3700 30144
rect 3752 30132 3758 30184
rect 4157 30175 4215 30181
rect 4157 30141 4169 30175
rect 4203 30141 4215 30175
rect 4157 30135 4215 30141
rect 4172 30104 4200 30135
rect 4246 30132 4252 30184
rect 4304 30172 4310 30184
rect 4525 30175 4583 30181
rect 4525 30172 4537 30175
rect 4304 30144 4537 30172
rect 4304 30132 4310 30144
rect 4525 30141 4537 30144
rect 4571 30141 4583 30175
rect 4525 30135 4583 30141
rect 7193 30175 7251 30181
rect 7193 30141 7205 30175
rect 7239 30172 7251 30175
rect 8202 30172 8208 30184
rect 7239 30144 8208 30172
rect 7239 30141 7251 30144
rect 7193 30135 7251 30141
rect 8202 30132 8208 30144
rect 8260 30172 8266 30184
rect 8757 30175 8815 30181
rect 8757 30172 8769 30175
rect 8260 30144 8769 30172
rect 8260 30132 8266 30144
rect 8757 30141 8769 30144
rect 8803 30141 8815 30175
rect 8757 30135 8815 30141
rect 9953 30175 10011 30181
rect 9953 30141 9965 30175
rect 9999 30141 10011 30175
rect 10134 30172 10140 30184
rect 10095 30144 10140 30172
rect 9953 30135 10011 30141
rect 3160 30076 4200 30104
rect 3160 30048 3188 30076
rect 5718 30064 5724 30116
rect 5776 30104 5782 30116
rect 7285 30107 7343 30113
rect 7285 30104 7297 30107
rect 5776 30076 7297 30104
rect 5776 30064 5782 30076
rect 7285 30073 7297 30076
rect 7331 30073 7343 30107
rect 9968 30104 9996 30135
rect 10134 30132 10140 30144
rect 10192 30132 10198 30184
rect 10594 30172 10600 30184
rect 10507 30144 10600 30172
rect 10594 30132 10600 30144
rect 10652 30132 10658 30184
rect 10781 30175 10839 30181
rect 10781 30141 10793 30175
rect 10827 30172 10839 30175
rect 10962 30172 10968 30184
rect 10827 30144 10968 30172
rect 10827 30141 10839 30144
rect 10781 30135 10839 30141
rect 10962 30132 10968 30144
rect 11020 30132 11026 30184
rect 11425 30175 11483 30181
rect 11425 30141 11437 30175
rect 11471 30172 11483 30175
rect 12434 30172 12440 30184
rect 11471 30144 12440 30172
rect 11471 30141 11483 30144
rect 11425 30135 11483 30141
rect 12434 30132 12440 30144
rect 12492 30132 12498 30184
rect 12986 30132 12992 30184
rect 13044 30172 13050 30184
rect 13081 30175 13139 30181
rect 13081 30172 13093 30175
rect 13044 30144 13093 30172
rect 13044 30132 13050 30144
rect 13081 30141 13093 30144
rect 13127 30141 13139 30175
rect 13081 30135 13139 30141
rect 13265 30175 13323 30181
rect 13265 30141 13277 30175
rect 13311 30172 13323 30175
rect 13740 30172 13768 30271
rect 14277 30243 14335 30249
rect 14277 30240 14289 30243
rect 13311 30144 13768 30172
rect 13832 30212 14289 30240
rect 13311 30141 13323 30144
rect 13265 30135 13323 30141
rect 10689 30107 10747 30113
rect 10689 30104 10701 30107
rect 9968 30076 10701 30104
rect 7285 30067 7343 30073
rect 10689 30073 10701 30076
rect 10735 30073 10747 30107
rect 10689 30067 10747 30073
rect 11606 30064 11612 30116
rect 11664 30104 11670 30116
rect 13832 30104 13860 30212
rect 14277 30209 14289 30212
rect 14323 30209 14335 30243
rect 14384 30240 14412 30280
rect 15105 30277 15117 30311
rect 15151 30308 15163 30311
rect 15286 30308 15292 30320
rect 15151 30280 15292 30308
rect 15151 30277 15163 30280
rect 15105 30271 15163 30277
rect 15286 30268 15292 30280
rect 15344 30268 15350 30320
rect 17402 30268 17408 30320
rect 17460 30308 17466 30320
rect 18233 30311 18291 30317
rect 18233 30308 18245 30311
rect 17460 30280 18245 30308
rect 17460 30268 17466 30280
rect 18233 30277 18245 30280
rect 18279 30277 18291 30311
rect 18233 30271 18291 30277
rect 15197 30243 15255 30249
rect 15197 30240 15209 30243
rect 14384 30212 15209 30240
rect 14277 30203 14335 30209
rect 15197 30209 15209 30212
rect 15243 30209 15255 30243
rect 15197 30203 15255 30209
rect 17954 30200 17960 30252
rect 18012 30240 18018 30252
rect 18693 30243 18751 30249
rect 18693 30240 18705 30243
rect 18012 30212 18705 30240
rect 18012 30200 18018 30212
rect 18693 30209 18705 30212
rect 18739 30209 18751 30243
rect 18693 30203 18751 30209
rect 18877 30243 18935 30249
rect 18877 30209 18889 30243
rect 18923 30240 18935 30243
rect 19150 30240 19156 30252
rect 18923 30212 19156 30240
rect 18923 30209 18935 30212
rect 18877 30203 18935 30209
rect 19150 30200 19156 30212
rect 19208 30240 19214 30252
rect 20346 30240 20352 30252
rect 19208 30212 20352 30240
rect 19208 30200 19214 30212
rect 20346 30200 20352 30212
rect 20404 30200 20410 30252
rect 21082 30240 21088 30252
rect 21043 30212 21088 30240
rect 21082 30200 21088 30212
rect 21140 30200 21146 30252
rect 22664 30249 22692 30348
rect 23566 30336 23572 30348
rect 23624 30336 23630 30388
rect 23934 30336 23940 30388
rect 23992 30376 23998 30388
rect 24443 30379 24501 30385
rect 24443 30376 24455 30379
rect 23992 30348 24455 30376
rect 23992 30336 23998 30348
rect 24443 30345 24455 30348
rect 24489 30376 24501 30379
rect 24762 30376 24768 30388
rect 24489 30348 24768 30376
rect 24489 30345 24501 30348
rect 24443 30339 24501 30345
rect 24762 30336 24768 30348
rect 24820 30336 24826 30388
rect 26053 30311 26111 30317
rect 26053 30277 26065 30311
rect 26099 30308 26111 30311
rect 27338 30308 27344 30320
rect 26099 30280 27344 30308
rect 26099 30277 26111 30280
rect 26053 30271 26111 30277
rect 27338 30268 27344 30280
rect 27396 30268 27402 30320
rect 22649 30243 22707 30249
rect 22649 30209 22661 30243
rect 22695 30209 22707 30243
rect 22649 30203 22707 30209
rect 23017 30243 23075 30249
rect 23017 30209 23029 30243
rect 23063 30240 23075 30243
rect 23474 30240 23480 30252
rect 23063 30212 23480 30240
rect 23063 30209 23075 30212
rect 23017 30203 23075 30209
rect 14182 30172 14188 30184
rect 14143 30144 14188 30172
rect 14182 30132 14188 30144
rect 14240 30132 14246 30184
rect 14918 30172 14924 30184
rect 14879 30144 14924 30172
rect 14918 30132 14924 30144
rect 14976 30132 14982 30184
rect 15013 30175 15071 30181
rect 15013 30141 15025 30175
rect 15059 30141 15071 30175
rect 18598 30172 18604 30184
rect 18559 30144 18604 30172
rect 15013 30135 15071 30141
rect 11664 30076 13860 30104
rect 11664 30064 11670 30076
rect 13906 30064 13912 30116
rect 13964 30104 13970 30116
rect 14093 30107 14151 30113
rect 14093 30104 14105 30107
rect 13964 30076 14105 30104
rect 13964 30064 13970 30076
rect 14093 30073 14105 30076
rect 14139 30073 14151 30107
rect 14093 30067 14151 30073
rect 2777 30039 2835 30045
rect 2777 30005 2789 30039
rect 2823 30036 2835 30039
rect 3142 30036 3148 30048
rect 2823 30008 3148 30036
rect 2823 30005 2835 30008
rect 2777 29999 2835 30005
rect 3142 29996 3148 30008
rect 3200 29996 3206 30048
rect 8570 29996 8576 30048
rect 8628 30036 8634 30048
rect 8849 30039 8907 30045
rect 8849 30036 8861 30039
rect 8628 30008 8861 30036
rect 8628 29996 8634 30008
rect 8849 30005 8861 30008
rect 8895 30005 8907 30039
rect 8849 29999 8907 30005
rect 10870 29996 10876 30048
rect 10928 30036 10934 30048
rect 11241 30039 11299 30045
rect 11241 30036 11253 30039
rect 10928 30008 11253 30036
rect 10928 29996 10934 30008
rect 11241 30005 11253 30008
rect 11287 30005 11299 30039
rect 11241 29999 11299 30005
rect 12802 29996 12808 30048
rect 12860 30036 12866 30048
rect 12986 30036 12992 30048
rect 12860 30008 12992 30036
rect 12860 29996 12866 30008
rect 12986 29996 12992 30008
rect 13044 30036 13050 30048
rect 15028 30036 15056 30135
rect 18598 30132 18604 30144
rect 18656 30132 18662 30184
rect 20990 30132 20996 30184
rect 21048 30172 21054 30184
rect 21358 30172 21364 30184
rect 21048 30144 21364 30172
rect 21048 30132 21054 30144
rect 21358 30132 21364 30144
rect 21416 30172 21422 30184
rect 21453 30175 21511 30181
rect 21453 30172 21465 30175
rect 21416 30144 21465 30172
rect 21416 30132 21422 30144
rect 21453 30141 21465 30144
rect 21499 30172 21511 30175
rect 22664 30172 22692 30203
rect 23474 30200 23480 30212
rect 23532 30200 23538 30252
rect 26602 30240 26608 30252
rect 26563 30212 26608 30240
rect 26602 30200 26608 30212
rect 26660 30200 26666 30252
rect 28350 30200 28356 30252
rect 28408 30240 28414 30252
rect 29365 30243 29423 30249
rect 29365 30240 29377 30243
rect 28408 30212 29377 30240
rect 28408 30200 28414 30212
rect 29365 30209 29377 30212
rect 29411 30209 29423 30243
rect 29914 30240 29920 30252
rect 29365 30203 29423 30209
rect 29840 30212 29920 30240
rect 21499 30144 22692 30172
rect 21499 30141 21511 30144
rect 21453 30135 21511 30141
rect 24854 30132 24860 30184
rect 24912 30172 24918 30184
rect 25317 30175 25375 30181
rect 25317 30172 25329 30175
rect 24912 30144 25329 30172
rect 24912 30132 24918 30144
rect 25317 30141 25329 30144
rect 25363 30172 25375 30175
rect 26142 30172 26148 30184
rect 25363 30144 26148 30172
rect 25363 30141 25375 30144
rect 25317 30135 25375 30141
rect 26142 30132 26148 30144
rect 26200 30132 26206 30184
rect 26234 30132 26240 30184
rect 26292 30172 26298 30184
rect 26513 30175 26571 30181
rect 26513 30172 26525 30175
rect 26292 30144 26525 30172
rect 26292 30132 26298 30144
rect 26513 30141 26525 30144
rect 26559 30141 26571 30175
rect 26513 30135 26571 30141
rect 29181 30175 29239 30181
rect 29181 30141 29193 30175
rect 29227 30172 29239 30175
rect 29546 30172 29552 30184
rect 29227 30144 29552 30172
rect 29227 30141 29239 30144
rect 29181 30135 29239 30141
rect 29546 30132 29552 30144
rect 29604 30132 29610 30184
rect 29840 30181 29868 30212
rect 29914 30200 29920 30212
rect 29972 30200 29978 30252
rect 29825 30175 29883 30181
rect 29825 30141 29837 30175
rect 29871 30141 29883 30175
rect 30006 30172 30012 30184
rect 29967 30144 30012 30172
rect 29825 30135 29883 30141
rect 30006 30132 30012 30144
rect 30064 30132 30070 30184
rect 24302 30104 24308 30116
rect 13044 30008 15056 30036
rect 13044 29996 13050 30008
rect 19610 29996 19616 30048
rect 19668 30045 19674 30048
rect 19668 30039 19717 30045
rect 19668 30005 19671 30039
rect 19705 30005 19717 30039
rect 20732 30036 20760 30090
rect 24058 30076 24308 30104
rect 24302 30064 24308 30076
rect 24360 30064 24366 30116
rect 21174 30036 21180 30048
rect 20732 30008 21180 30036
rect 19668 29999 19717 30005
rect 19668 29996 19674 29999
rect 21174 29996 21180 30008
rect 21232 29996 21238 30048
rect 25501 30039 25559 30045
rect 25501 30005 25513 30039
rect 25547 30036 25559 30039
rect 25866 30036 25872 30048
rect 25547 30008 25872 30036
rect 25547 30005 25559 30008
rect 25501 29999 25559 30005
rect 25866 29996 25872 30008
rect 25924 29996 25930 30048
rect 26418 30036 26424 30048
rect 26379 30008 26424 30036
rect 26418 29996 26424 30008
rect 26476 29996 26482 30048
rect 1104 29946 34316 29968
rect 1104 29894 12052 29946
rect 12104 29894 12116 29946
rect 12168 29894 12180 29946
rect 12232 29894 12244 29946
rect 12296 29894 23123 29946
rect 23175 29894 23187 29946
rect 23239 29894 23251 29946
rect 23303 29894 23315 29946
rect 23367 29894 34316 29946
rect 1104 29872 34316 29894
rect 2961 29835 3019 29841
rect 2961 29801 2973 29835
rect 3007 29832 3019 29835
rect 3234 29832 3240 29844
rect 3007 29804 3240 29832
rect 3007 29801 3019 29804
rect 2961 29795 3019 29801
rect 3234 29792 3240 29804
rect 3292 29792 3298 29844
rect 5626 29832 5632 29844
rect 5587 29804 5632 29832
rect 5626 29792 5632 29804
rect 5684 29792 5690 29844
rect 9766 29832 9772 29844
rect 9727 29804 9772 29832
rect 9766 29792 9772 29804
rect 9824 29792 9830 29844
rect 10962 29832 10968 29844
rect 10923 29804 10968 29832
rect 10962 29792 10968 29804
rect 11020 29792 11026 29844
rect 12621 29835 12679 29841
rect 12621 29801 12633 29835
rect 12667 29832 12679 29835
rect 13078 29832 13084 29844
rect 12667 29804 13084 29832
rect 12667 29801 12679 29804
rect 12621 29795 12679 29801
rect 13078 29792 13084 29804
rect 13136 29792 13142 29844
rect 14921 29835 14979 29841
rect 14921 29801 14933 29835
rect 14967 29832 14979 29835
rect 16114 29832 16120 29844
rect 14967 29804 16120 29832
rect 14967 29801 14979 29804
rect 14921 29795 14979 29801
rect 16114 29792 16120 29804
rect 16172 29792 16178 29844
rect 21174 29832 21180 29844
rect 18616 29804 21180 29832
rect 4709 29767 4767 29773
rect 4709 29764 4721 29767
rect 3160 29736 4721 29764
rect 3160 29708 3188 29736
rect 4709 29733 4721 29736
rect 4755 29733 4767 29767
rect 11333 29767 11391 29773
rect 4709 29727 4767 29733
rect 5552 29736 11284 29764
rect 3142 29696 3148 29708
rect 3103 29668 3148 29696
rect 3142 29656 3148 29668
rect 3200 29656 3206 29708
rect 4617 29699 4675 29705
rect 4617 29665 4629 29699
rect 4663 29696 4675 29699
rect 5552 29696 5580 29736
rect 5718 29696 5724 29708
rect 4663 29668 5580 29696
rect 5679 29668 5724 29696
rect 4663 29665 4675 29668
rect 4617 29659 4675 29665
rect 5718 29656 5724 29668
rect 5776 29656 5782 29708
rect 5902 29696 5908 29708
rect 5863 29668 5908 29696
rect 5902 29656 5908 29668
rect 5960 29656 5966 29708
rect 7745 29699 7803 29705
rect 7745 29665 7757 29699
rect 7791 29696 7803 29699
rect 8018 29696 8024 29708
rect 7791 29668 8024 29696
rect 7791 29665 7803 29668
rect 7745 29659 7803 29665
rect 8018 29656 8024 29668
rect 8076 29656 8082 29708
rect 8570 29656 8576 29708
rect 8628 29696 8634 29708
rect 9493 29699 9551 29705
rect 9493 29696 9505 29699
rect 8628 29668 9505 29696
rect 8628 29656 8634 29668
rect 9493 29665 9505 29668
rect 9539 29665 9551 29699
rect 10226 29696 10232 29708
rect 10187 29668 10232 29696
rect 9493 29659 9551 29665
rect 10226 29656 10232 29668
rect 10284 29656 10290 29708
rect 10413 29699 10471 29705
rect 10413 29665 10425 29699
rect 10459 29696 10471 29699
rect 10594 29696 10600 29708
rect 10459 29668 10600 29696
rect 10459 29665 10471 29668
rect 10413 29659 10471 29665
rect 3329 29631 3387 29637
rect 3329 29597 3341 29631
rect 3375 29628 3387 29631
rect 4338 29628 4344 29640
rect 3375 29600 4344 29628
rect 3375 29597 3387 29600
rect 3329 29591 3387 29597
rect 4338 29588 4344 29600
rect 4396 29588 4402 29640
rect 4893 29631 4951 29637
rect 4893 29597 4905 29631
rect 4939 29628 4951 29631
rect 4982 29628 4988 29640
rect 4939 29600 4988 29628
rect 4939 29597 4951 29600
rect 4893 29591 4951 29597
rect 4982 29588 4988 29600
rect 5040 29588 5046 29640
rect 7469 29631 7527 29637
rect 7469 29597 7481 29631
rect 7515 29597 7527 29631
rect 7650 29628 7656 29640
rect 7611 29600 7656 29628
rect 7469 29591 7527 29597
rect 7484 29560 7512 29591
rect 7650 29588 7656 29600
rect 7708 29588 7714 29640
rect 9769 29631 9827 29637
rect 9769 29597 9781 29631
rect 9815 29628 9827 29631
rect 10321 29631 10379 29637
rect 10321 29628 10333 29631
rect 9815 29600 10333 29628
rect 9815 29597 9827 29600
rect 9769 29591 9827 29597
rect 10321 29597 10333 29600
rect 10367 29597 10379 29631
rect 10321 29591 10379 29597
rect 9585 29563 9643 29569
rect 7484 29532 9444 29560
rect 3418 29452 3424 29504
rect 3476 29492 3482 29504
rect 4249 29495 4307 29501
rect 4249 29492 4261 29495
rect 3476 29464 4261 29492
rect 3476 29452 3482 29464
rect 4249 29461 4261 29464
rect 4295 29461 4307 29495
rect 4249 29455 4307 29461
rect 8113 29495 8171 29501
rect 8113 29461 8125 29495
rect 8159 29492 8171 29495
rect 9122 29492 9128 29504
rect 8159 29464 9128 29492
rect 8159 29461 8171 29464
rect 8113 29455 8171 29461
rect 9122 29452 9128 29464
rect 9180 29452 9186 29504
rect 9416 29492 9444 29532
rect 9585 29529 9597 29563
rect 9631 29560 9643 29563
rect 9858 29560 9864 29572
rect 9631 29532 9864 29560
rect 9631 29529 9643 29532
rect 9585 29523 9643 29529
rect 9858 29520 9864 29532
rect 9916 29560 9922 29572
rect 10428 29560 10456 29659
rect 10594 29656 10600 29668
rect 10652 29656 10658 29708
rect 11256 29696 11284 29736
rect 11333 29733 11345 29767
rect 11379 29764 11391 29767
rect 11422 29764 11428 29776
rect 11379 29736 11428 29764
rect 11379 29733 11391 29736
rect 11333 29727 11391 29733
rect 11422 29724 11428 29736
rect 11480 29724 11486 29776
rect 12529 29767 12587 29773
rect 12529 29733 12541 29767
rect 12575 29764 12587 29767
rect 12710 29764 12716 29776
rect 12575 29736 12716 29764
rect 12575 29733 12587 29736
rect 12529 29727 12587 29733
rect 12710 29724 12716 29736
rect 12768 29724 12774 29776
rect 16390 29724 16396 29776
rect 16448 29773 16454 29776
rect 16448 29764 16460 29773
rect 16758 29764 16764 29776
rect 16448 29736 16764 29764
rect 16448 29727 16460 29736
rect 16448 29724 16454 29727
rect 16758 29724 16764 29736
rect 16816 29724 16822 29776
rect 14366 29696 14372 29708
rect 11256 29668 12434 29696
rect 11425 29631 11483 29637
rect 11425 29597 11437 29631
rect 11471 29597 11483 29631
rect 11606 29628 11612 29640
rect 11567 29600 11612 29628
rect 11425 29591 11483 29597
rect 9916 29532 10456 29560
rect 11440 29560 11468 29591
rect 11606 29588 11612 29600
rect 11664 29588 11670 29640
rect 12406 29628 12434 29668
rect 12636 29668 14372 29696
rect 12636 29628 12664 29668
rect 14366 29656 14372 29668
rect 14424 29656 14430 29708
rect 14737 29699 14795 29705
rect 14737 29665 14749 29699
rect 14783 29665 14795 29699
rect 14737 29659 14795 29665
rect 12406 29600 12664 29628
rect 12805 29631 12863 29637
rect 12805 29597 12817 29631
rect 12851 29628 12863 29631
rect 12894 29628 12900 29640
rect 12851 29600 12900 29628
rect 12851 29597 12863 29600
rect 12805 29591 12863 29597
rect 12894 29588 12900 29600
rect 12952 29588 12958 29640
rect 12161 29563 12219 29569
rect 12161 29560 12173 29563
rect 11440 29532 12173 29560
rect 9916 29520 9922 29532
rect 12161 29529 12173 29532
rect 12207 29529 12219 29563
rect 12161 29523 12219 29529
rect 12434 29520 12440 29572
rect 12492 29560 12498 29572
rect 14752 29560 14780 29659
rect 16114 29656 16120 29708
rect 16172 29696 16178 29708
rect 16172 29668 16712 29696
rect 16172 29656 16178 29668
rect 16684 29637 16712 29668
rect 18414 29656 18420 29708
rect 18472 29696 18478 29708
rect 18616 29696 18644 29804
rect 21174 29792 21180 29804
rect 21232 29832 21238 29844
rect 21232 29804 21864 29832
rect 21232 29792 21238 29804
rect 21836 29750 21864 29804
rect 31754 29792 31760 29844
rect 31812 29792 31818 29844
rect 26418 29764 26424 29776
rect 26160 29736 26424 29764
rect 18472 29668 18644 29696
rect 18472 29656 18478 29668
rect 24762 29656 24768 29708
rect 24820 29696 24826 29708
rect 25225 29699 25283 29705
rect 25225 29696 25237 29699
rect 24820 29668 25237 29696
rect 24820 29656 24826 29668
rect 25225 29665 25237 29668
rect 25271 29665 25283 29699
rect 25225 29659 25283 29665
rect 25498 29656 25504 29708
rect 25556 29696 25562 29708
rect 26160 29705 26188 29736
rect 26418 29724 26424 29736
rect 26476 29724 26482 29776
rect 31772 29750 31800 29792
rect 26053 29699 26111 29705
rect 26053 29696 26065 29699
rect 25556 29668 26065 29696
rect 25556 29656 25562 29668
rect 26053 29665 26065 29668
rect 26099 29665 26111 29699
rect 26053 29659 26111 29665
rect 26145 29699 26203 29705
rect 26145 29665 26157 29699
rect 26191 29665 26203 29699
rect 26145 29659 26203 29665
rect 26234 29656 26240 29708
rect 26292 29696 26298 29708
rect 27985 29699 28043 29705
rect 27985 29696 27997 29699
rect 26292 29668 26337 29696
rect 27540 29668 27997 29696
rect 26292 29656 26298 29668
rect 16669 29631 16727 29637
rect 16669 29597 16681 29631
rect 16715 29628 16727 29631
rect 17218 29628 17224 29640
rect 16715 29600 17224 29628
rect 16715 29597 16727 29600
rect 16669 29591 16727 29597
rect 17218 29588 17224 29600
rect 17276 29588 17282 29640
rect 17589 29631 17647 29637
rect 17589 29597 17601 29631
rect 17635 29628 17647 29631
rect 18322 29628 18328 29640
rect 17635 29600 18328 29628
rect 17635 29597 17647 29600
rect 17589 29591 17647 29597
rect 18322 29588 18328 29600
rect 18380 29588 18386 29640
rect 18598 29588 18604 29640
rect 18656 29628 18662 29640
rect 19015 29631 19073 29637
rect 19015 29628 19027 29631
rect 18656 29600 19027 29628
rect 18656 29588 18662 29600
rect 19015 29597 19027 29600
rect 19061 29597 19073 29631
rect 19015 29591 19073 29597
rect 20898 29588 20904 29640
rect 20956 29628 20962 29640
rect 21085 29631 21143 29637
rect 21085 29628 21097 29631
rect 20956 29600 21097 29628
rect 20956 29588 20962 29600
rect 21085 29597 21097 29600
rect 21131 29597 21143 29631
rect 21450 29628 21456 29640
rect 21411 29600 21456 29628
rect 21085 29591 21143 29597
rect 21450 29588 21456 29600
rect 21508 29588 21514 29640
rect 12492 29532 14780 29560
rect 12492 29520 12498 29532
rect 24854 29520 24860 29572
rect 24912 29560 24918 29572
rect 25869 29563 25927 29569
rect 25869 29560 25881 29563
rect 24912 29532 25881 29560
rect 24912 29520 24918 29532
rect 25869 29529 25881 29532
rect 25915 29529 25927 29563
rect 25869 29523 25927 29529
rect 26234 29520 26240 29572
rect 26292 29560 26298 29572
rect 27540 29560 27568 29668
rect 27985 29665 27997 29668
rect 28031 29665 28043 29699
rect 28350 29696 28356 29708
rect 28311 29668 28356 29696
rect 27985 29659 28043 29665
rect 28350 29656 28356 29668
rect 28408 29656 28414 29708
rect 28813 29699 28871 29705
rect 28813 29665 28825 29699
rect 28859 29696 28871 29699
rect 28994 29696 29000 29708
rect 28859 29668 29000 29696
rect 28859 29665 28871 29668
rect 28813 29659 28871 29665
rect 28994 29656 29000 29668
rect 29052 29656 29058 29708
rect 27614 29588 27620 29640
rect 27672 29628 27678 29640
rect 30653 29631 30711 29637
rect 30653 29628 30665 29631
rect 27672 29600 30665 29628
rect 27672 29588 27678 29600
rect 30653 29597 30665 29600
rect 30699 29597 30711 29631
rect 30926 29628 30932 29640
rect 30887 29600 30932 29628
rect 30653 29591 30711 29597
rect 30926 29588 30932 29600
rect 30984 29588 30990 29640
rect 26292 29532 27568 29560
rect 26292 29520 26298 29532
rect 27890 29520 27896 29572
rect 27948 29560 27954 29572
rect 27948 29532 27993 29560
rect 27948 29520 27954 29532
rect 12894 29492 12900 29504
rect 9416 29464 12900 29492
rect 12894 29452 12900 29464
rect 12952 29492 12958 29504
rect 13722 29492 13728 29504
rect 12952 29464 13728 29492
rect 12952 29452 12958 29464
rect 13722 29452 13728 29464
rect 13780 29452 13786 29504
rect 15289 29495 15347 29501
rect 15289 29461 15301 29495
rect 15335 29492 15347 29495
rect 16666 29492 16672 29504
rect 15335 29464 16672 29492
rect 15335 29461 15347 29464
rect 15289 29455 15347 29461
rect 16666 29452 16672 29464
rect 16724 29452 16730 29504
rect 20530 29452 20536 29504
rect 20588 29492 20594 29504
rect 22002 29492 22008 29504
rect 20588 29464 22008 29492
rect 20588 29452 20594 29464
rect 22002 29452 22008 29464
rect 22060 29492 22066 29504
rect 22879 29495 22937 29501
rect 22879 29492 22891 29495
rect 22060 29464 22891 29492
rect 22060 29452 22066 29464
rect 22879 29461 22891 29464
rect 22925 29461 22937 29495
rect 22879 29455 22937 29461
rect 25130 29452 25136 29504
rect 25188 29492 25194 29504
rect 25317 29495 25375 29501
rect 25317 29492 25329 29495
rect 25188 29464 25329 29492
rect 25188 29452 25194 29464
rect 25317 29461 25329 29464
rect 25363 29461 25375 29495
rect 25317 29455 25375 29461
rect 31294 29452 31300 29504
rect 31352 29492 31358 29504
rect 32401 29495 32459 29501
rect 32401 29492 32413 29495
rect 31352 29464 32413 29492
rect 31352 29452 31358 29464
rect 32401 29461 32413 29464
rect 32447 29461 32459 29495
rect 32401 29455 32459 29461
rect 1104 29402 34316 29424
rect 1104 29350 6517 29402
rect 6569 29350 6581 29402
rect 6633 29350 6645 29402
rect 6697 29350 6709 29402
rect 6761 29350 17588 29402
rect 17640 29350 17652 29402
rect 17704 29350 17716 29402
rect 17768 29350 17780 29402
rect 17832 29350 28658 29402
rect 28710 29350 28722 29402
rect 28774 29350 28786 29402
rect 28838 29350 28850 29402
rect 28902 29350 34316 29402
rect 1104 29328 34316 29350
rect 1949 29291 2007 29297
rect 1949 29257 1961 29291
rect 1995 29288 2007 29291
rect 8018 29288 8024 29300
rect 1995 29260 7604 29288
rect 7979 29260 8024 29288
rect 1995 29257 2007 29260
rect 1949 29251 2007 29257
rect 4062 29220 4068 29232
rect 3252 29192 4068 29220
rect 3252 29164 3280 29192
rect 4062 29180 4068 29192
rect 4120 29180 4126 29232
rect 5442 29180 5448 29232
rect 5500 29220 5506 29232
rect 5537 29223 5595 29229
rect 5537 29220 5549 29223
rect 5500 29192 5549 29220
rect 5500 29180 5506 29192
rect 5537 29189 5549 29192
rect 5583 29189 5595 29223
rect 5537 29183 5595 29189
rect 3234 29152 3240 29164
rect 3195 29124 3240 29152
rect 3234 29112 3240 29124
rect 3292 29112 3298 29164
rect 3418 29152 3424 29164
rect 3379 29124 3424 29152
rect 3418 29112 3424 29124
rect 3476 29112 3482 29164
rect 7190 29112 7196 29164
rect 7248 29152 7254 29164
rect 7576 29161 7604 29260
rect 8018 29248 8024 29260
rect 8076 29248 8082 29300
rect 9858 29288 9864 29300
rect 9819 29260 9864 29288
rect 9858 29248 9864 29260
rect 9916 29248 9922 29300
rect 12434 29248 12440 29300
rect 12492 29288 12498 29300
rect 12710 29288 12716 29300
rect 12492 29260 12537 29288
rect 12671 29260 12716 29288
rect 12492 29248 12498 29260
rect 12710 29248 12716 29260
rect 12768 29248 12774 29300
rect 18322 29288 18328 29300
rect 18283 29260 18328 29288
rect 18322 29248 18328 29260
rect 18380 29248 18386 29300
rect 20898 29248 20904 29300
rect 20956 29288 20962 29300
rect 23385 29291 23443 29297
rect 23385 29288 23397 29291
rect 20956 29260 23397 29288
rect 20956 29248 20962 29260
rect 23385 29257 23397 29260
rect 23431 29257 23443 29291
rect 25314 29288 25320 29300
rect 25275 29260 25320 29288
rect 23385 29251 23443 29257
rect 25314 29248 25320 29260
rect 25372 29248 25378 29300
rect 25498 29288 25504 29300
rect 25459 29260 25504 29288
rect 25498 29248 25504 29260
rect 25556 29248 25562 29300
rect 30653 29291 30711 29297
rect 30653 29257 30665 29291
rect 30699 29288 30711 29291
rect 30926 29288 30932 29300
rect 30699 29260 30932 29288
rect 30699 29257 30711 29260
rect 30653 29251 30711 29257
rect 30926 29248 30932 29260
rect 30984 29248 30990 29300
rect 7650 29180 7656 29232
rect 7708 29220 7714 29232
rect 8481 29223 8539 29229
rect 8481 29220 8493 29223
rect 7708 29192 8493 29220
rect 7708 29180 7714 29192
rect 8481 29189 8493 29192
rect 8527 29189 8539 29223
rect 11882 29220 11888 29232
rect 8481 29183 8539 29189
rect 9140 29192 11888 29220
rect 7377 29155 7435 29161
rect 7377 29152 7389 29155
rect 7248 29124 7389 29152
rect 7248 29112 7254 29124
rect 7377 29121 7389 29124
rect 7423 29121 7435 29155
rect 7377 29115 7435 29121
rect 7561 29155 7619 29161
rect 7561 29121 7573 29155
rect 7607 29121 7619 29155
rect 7561 29115 7619 29121
rect 8202 29112 8208 29164
rect 8260 29152 8266 29164
rect 9140 29161 9168 29192
rect 11882 29180 11888 29192
rect 11940 29220 11946 29232
rect 12526 29220 12532 29232
rect 11940 29192 12532 29220
rect 11940 29180 11946 29192
rect 12526 29180 12532 29192
rect 12584 29220 12590 29232
rect 26513 29223 26571 29229
rect 12584 29192 14412 29220
rect 12584 29180 12590 29192
rect 8941 29155 8999 29161
rect 8941 29152 8953 29155
rect 8260 29124 8953 29152
rect 8260 29112 8266 29124
rect 8941 29121 8953 29124
rect 8987 29121 8999 29155
rect 8941 29115 8999 29121
rect 9125 29155 9183 29161
rect 9125 29121 9137 29155
rect 9171 29121 9183 29155
rect 9125 29115 9183 29121
rect 13170 29112 13176 29164
rect 13228 29152 13234 29164
rect 14384 29161 14412 29192
rect 26513 29189 26525 29223
rect 26559 29220 26571 29223
rect 27614 29220 27620 29232
rect 26559 29192 27620 29220
rect 26559 29189 26571 29192
rect 26513 29183 26571 29189
rect 27614 29180 27620 29192
rect 27672 29220 27678 29232
rect 27672 29192 28028 29220
rect 27672 29180 27678 29192
rect 13265 29155 13323 29161
rect 13265 29152 13277 29155
rect 13228 29124 13277 29152
rect 13228 29112 13234 29124
rect 13265 29121 13277 29124
rect 13311 29121 13323 29155
rect 13265 29115 13323 29121
rect 14369 29155 14427 29161
rect 14369 29121 14381 29155
rect 14415 29121 14427 29155
rect 14369 29115 14427 29121
rect 16666 29112 16672 29164
rect 16724 29152 16730 29164
rect 16724 29124 17540 29152
rect 16724 29112 16730 29124
rect 1762 29084 1768 29096
rect 1723 29056 1768 29084
rect 1762 29044 1768 29056
rect 1820 29044 1826 29096
rect 3050 29044 3056 29096
rect 3108 29084 3114 29096
rect 3326 29084 3332 29096
rect 3108 29056 3332 29084
rect 3108 29044 3114 29056
rect 3326 29044 3332 29056
rect 3384 29044 3390 29096
rect 3513 29087 3571 29093
rect 3513 29053 3525 29087
rect 3559 29084 3571 29087
rect 4065 29087 4123 29093
rect 4065 29084 4077 29087
rect 3559 29056 4077 29084
rect 3559 29053 3571 29056
rect 3513 29047 3571 29053
rect 4065 29053 4077 29056
rect 4111 29053 4123 29087
rect 4246 29084 4252 29096
rect 4207 29056 4252 29084
rect 4065 29047 4123 29053
rect 4246 29044 4252 29056
rect 4304 29044 4310 29096
rect 4338 29044 4344 29096
rect 4396 29084 4402 29096
rect 5261 29087 5319 29093
rect 4396 29056 4441 29084
rect 4396 29044 4402 29056
rect 5261 29053 5273 29087
rect 5307 29053 5319 29087
rect 5261 29047 5319 29053
rect 5353 29087 5411 29093
rect 5353 29053 5365 29087
rect 5399 29053 5411 29087
rect 5353 29047 5411 29053
rect 5629 29087 5687 29093
rect 5629 29053 5641 29087
rect 5675 29084 5687 29087
rect 5718 29084 5724 29096
rect 5675 29056 5724 29084
rect 5675 29053 5687 29056
rect 5629 29047 5687 29053
rect 3050 28948 3056 28960
rect 3011 28920 3056 28948
rect 3050 28908 3056 28920
rect 3108 28908 3114 28960
rect 5074 28948 5080 28960
rect 5035 28920 5080 28948
rect 5074 28908 5080 28920
rect 5132 28908 5138 28960
rect 5276 28948 5304 29047
rect 5368 29016 5396 29047
rect 5718 29044 5724 29056
rect 5776 29044 5782 29096
rect 7650 29084 7656 29096
rect 7611 29056 7656 29084
rect 7650 29044 7656 29056
rect 7708 29044 7714 29096
rect 9490 29044 9496 29096
rect 9548 29084 9554 29096
rect 9769 29087 9827 29093
rect 9769 29084 9781 29087
rect 9548 29056 9781 29084
rect 9548 29044 9554 29056
rect 9769 29053 9781 29056
rect 9815 29053 9827 29087
rect 9769 29047 9827 29053
rect 9950 29044 9956 29096
rect 10008 29084 10014 29096
rect 10505 29087 10563 29093
rect 10505 29084 10517 29087
rect 10008 29056 10517 29084
rect 10008 29044 10014 29056
rect 10505 29053 10517 29056
rect 10551 29053 10563 29087
rect 10686 29084 10692 29096
rect 10647 29056 10692 29084
rect 10505 29047 10563 29053
rect 10686 29044 10692 29056
rect 10744 29044 10750 29096
rect 12621 29087 12679 29093
rect 12621 29053 12633 29087
rect 12667 29084 12679 29087
rect 12894 29084 12900 29096
rect 12667 29056 12900 29084
rect 12667 29053 12679 29056
rect 12621 29047 12679 29053
rect 12894 29044 12900 29056
rect 12952 29044 12958 29096
rect 13078 29084 13084 29096
rect 13039 29056 13084 29084
rect 13078 29044 13084 29056
rect 13136 29044 13142 29096
rect 16758 29044 16764 29096
rect 16816 29084 16822 29096
rect 17512 29093 17540 29124
rect 18598 29112 18604 29164
rect 18656 29152 18662 29164
rect 18785 29155 18843 29161
rect 18785 29152 18797 29155
rect 18656 29124 18797 29152
rect 18656 29112 18662 29124
rect 18785 29121 18797 29124
rect 18831 29121 18843 29155
rect 18785 29115 18843 29121
rect 18969 29155 19027 29161
rect 18969 29121 18981 29155
rect 19015 29152 19027 29155
rect 19150 29152 19156 29164
rect 19015 29124 19156 29152
rect 19015 29121 19027 29124
rect 18969 29115 19027 29121
rect 19150 29112 19156 29124
rect 19208 29112 19214 29164
rect 24578 29152 24584 29164
rect 23584 29124 24584 29152
rect 17313 29087 17371 29093
rect 17313 29084 17325 29087
rect 16816 29056 17325 29084
rect 16816 29044 16822 29056
rect 17313 29053 17325 29056
rect 17359 29053 17371 29087
rect 17313 29047 17371 29053
rect 17497 29087 17555 29093
rect 17497 29053 17509 29087
rect 17543 29053 17555 29087
rect 17497 29047 17555 29053
rect 18693 29087 18751 29093
rect 18693 29053 18705 29087
rect 18739 29084 18751 29087
rect 19610 29084 19616 29096
rect 18739 29056 19616 29084
rect 18739 29053 18751 29056
rect 18693 29047 18751 29053
rect 19610 29044 19616 29056
rect 19668 29044 19674 29096
rect 20349 29087 20407 29093
rect 20349 29053 20361 29087
rect 20395 29084 20407 29087
rect 20438 29084 20444 29096
rect 20395 29056 20444 29084
rect 20395 29053 20407 29056
rect 20349 29047 20407 29053
rect 20438 29044 20444 29056
rect 20496 29044 20502 29096
rect 20530 29044 20536 29096
rect 20588 29084 20594 29096
rect 23584 29093 23612 29124
rect 24578 29112 24584 29124
rect 24636 29152 24642 29164
rect 28000 29161 28028 29192
rect 32398 29180 32404 29232
rect 32456 29220 32462 29232
rect 33413 29223 33471 29229
rect 33413 29220 33425 29223
rect 32456 29192 33425 29220
rect 32456 29180 32462 29192
rect 33413 29189 33425 29192
rect 33459 29189 33471 29223
rect 33413 29183 33471 29189
rect 27985 29155 28043 29161
rect 24636 29124 26372 29152
rect 24636 29112 24642 29124
rect 26344 29093 26372 29124
rect 27985 29121 27997 29155
rect 28031 29121 28043 29155
rect 31202 29152 31208 29164
rect 31163 29124 31208 29152
rect 27985 29115 28043 29121
rect 31202 29112 31208 29124
rect 31260 29112 31266 29164
rect 23569 29087 23627 29093
rect 20588 29056 20633 29084
rect 20588 29044 20594 29056
rect 23569 29053 23581 29087
rect 23615 29053 23627 29087
rect 23569 29047 23627 29053
rect 24213 29087 24271 29093
rect 24213 29053 24225 29087
rect 24259 29053 24271 29087
rect 24213 29047 24271 29053
rect 24397 29087 24455 29093
rect 24397 29053 24409 29087
rect 24443 29053 24455 29087
rect 24397 29047 24455 29053
rect 26329 29087 26387 29093
rect 26329 29053 26341 29087
rect 26375 29053 26387 29087
rect 26329 29047 26387 29053
rect 5534 29016 5540 29028
rect 5368 28988 5540 29016
rect 5534 28976 5540 28988
rect 5592 28976 5598 29028
rect 6822 29016 6828 29028
rect 5644 28988 6828 29016
rect 5644 28948 5672 28988
rect 6822 28976 6828 28988
rect 6880 28976 6886 29028
rect 12710 28976 12716 29028
rect 12768 29016 12774 29028
rect 13173 29019 13231 29025
rect 13173 29016 13185 29019
rect 12768 28988 13185 29016
rect 12768 28976 12774 28988
rect 13173 28985 13185 28988
rect 13219 28985 13231 29019
rect 13173 28979 13231 28985
rect 17402 28976 17408 29028
rect 17460 29016 17466 29028
rect 17681 29019 17739 29025
rect 17681 29016 17693 29019
rect 17460 28988 17693 29016
rect 17460 28976 17466 28988
rect 17681 28985 17693 28988
rect 17727 28985 17739 29019
rect 17681 28979 17739 28985
rect 22554 28976 22560 29028
rect 22612 29016 22618 29028
rect 24228 29016 24256 29047
rect 22612 28988 24256 29016
rect 24412 29016 24440 29047
rect 29362 29044 29368 29096
rect 29420 29084 29426 29096
rect 30098 29084 30104 29096
rect 29420 29056 30104 29084
rect 29420 29044 29426 29056
rect 30098 29044 30104 29056
rect 30156 29044 30162 29096
rect 31021 29087 31079 29093
rect 31021 29053 31033 29087
rect 31067 29084 31079 29087
rect 31294 29084 31300 29096
rect 31067 29056 31300 29084
rect 31067 29053 31079 29056
rect 31021 29047 31079 29053
rect 31294 29044 31300 29056
rect 31352 29044 31358 29096
rect 33594 29084 33600 29096
rect 33555 29056 33600 29084
rect 33594 29044 33600 29056
rect 33652 29044 33658 29096
rect 25130 29016 25136 29028
rect 24412 28988 25136 29016
rect 22612 28976 22618 28988
rect 25130 28976 25136 28988
rect 25188 28976 25194 29028
rect 28258 29016 28264 29028
rect 28219 28988 28264 29016
rect 28258 28976 28264 28988
rect 28316 28976 28322 29028
rect 30282 29016 30288 29028
rect 29748 28988 30288 29016
rect 8846 28948 8852 28960
rect 5276 28920 5672 28948
rect 8807 28920 8852 28948
rect 8846 28908 8852 28920
rect 8904 28908 8910 28960
rect 10597 28951 10655 28957
rect 10597 28917 10609 28951
rect 10643 28948 10655 28951
rect 10962 28948 10968 28960
rect 10643 28920 10968 28948
rect 10643 28917 10655 28920
rect 10597 28911 10655 28917
rect 10962 28908 10968 28920
rect 11020 28908 11026 28960
rect 14550 28948 14556 28960
rect 14511 28920 14556 28948
rect 14550 28908 14556 28920
rect 14608 28908 14614 28960
rect 14642 28908 14648 28960
rect 14700 28948 14706 28960
rect 15010 28948 15016 28960
rect 14700 28920 14745 28948
rect 14971 28920 15016 28948
rect 14700 28908 14706 28920
rect 15010 28908 15016 28920
rect 15068 28908 15074 28960
rect 20346 28948 20352 28960
rect 20307 28920 20352 28948
rect 20346 28908 20352 28920
rect 20404 28908 20410 28960
rect 24302 28948 24308 28960
rect 24263 28920 24308 28948
rect 24302 28908 24308 28920
rect 24360 28908 24366 28960
rect 25338 28951 25396 28957
rect 25338 28917 25350 28951
rect 25384 28948 25396 28951
rect 25590 28948 25596 28960
rect 25384 28920 25596 28948
rect 25384 28917 25396 28920
rect 25338 28911 25396 28917
rect 25590 28908 25596 28920
rect 25648 28908 25654 28960
rect 29748 28957 29776 28988
rect 30282 28976 30288 28988
rect 30340 29016 30346 29028
rect 31113 29019 31171 29025
rect 31113 29016 31125 29019
rect 30340 28988 31125 29016
rect 30340 28976 30346 28988
rect 31113 28985 31125 28988
rect 31159 28985 31171 29019
rect 31113 28979 31171 28985
rect 29733 28951 29791 28957
rect 29733 28917 29745 28951
rect 29779 28917 29791 28951
rect 29733 28911 29791 28917
rect 1104 28858 34316 28880
rect 1104 28806 12052 28858
rect 12104 28806 12116 28858
rect 12168 28806 12180 28858
rect 12232 28806 12244 28858
rect 12296 28806 23123 28858
rect 23175 28806 23187 28858
rect 23239 28806 23251 28858
rect 23303 28806 23315 28858
rect 23367 28806 34316 28858
rect 1104 28784 34316 28806
rect 3145 28747 3203 28753
rect 3145 28713 3157 28747
rect 3191 28744 3203 28747
rect 4246 28744 4252 28756
rect 3191 28716 4252 28744
rect 3191 28713 3203 28716
rect 3145 28707 3203 28713
rect 4246 28704 4252 28716
rect 4304 28704 4310 28756
rect 5718 28704 5724 28756
rect 5776 28744 5782 28756
rect 6181 28747 6239 28753
rect 6181 28744 6193 28747
rect 5776 28716 6193 28744
rect 5776 28704 5782 28716
rect 6181 28713 6193 28716
rect 6227 28713 6239 28747
rect 6181 28707 6239 28713
rect 8573 28747 8631 28753
rect 8573 28713 8585 28747
rect 8619 28744 8631 28747
rect 8846 28744 8852 28756
rect 8619 28716 8852 28744
rect 8619 28713 8631 28716
rect 8573 28707 8631 28713
rect 8846 28704 8852 28716
rect 8904 28704 8910 28756
rect 9122 28704 9128 28756
rect 9180 28744 9186 28756
rect 9769 28747 9827 28753
rect 9769 28744 9781 28747
rect 9180 28716 9781 28744
rect 9180 28704 9186 28716
rect 9769 28713 9781 28716
rect 9815 28713 9827 28747
rect 10226 28744 10232 28756
rect 10187 28716 10232 28744
rect 9769 28707 9827 28713
rect 10226 28704 10232 28716
rect 10284 28704 10290 28756
rect 12345 28747 12403 28753
rect 12345 28713 12357 28747
rect 12391 28744 12403 28747
rect 14550 28744 14556 28756
rect 12391 28716 14556 28744
rect 12391 28713 12403 28716
rect 12345 28707 12403 28713
rect 2032 28679 2090 28685
rect 2032 28645 2044 28679
rect 2078 28676 2090 28679
rect 3050 28676 3056 28688
rect 2078 28648 3056 28676
rect 2078 28645 2090 28648
rect 2032 28639 2090 28645
rect 3050 28636 3056 28648
rect 3108 28636 3114 28688
rect 5074 28685 5080 28688
rect 5068 28676 5080 28685
rect 5035 28648 5080 28676
rect 5068 28639 5080 28648
rect 5074 28636 5080 28639
rect 5132 28636 5138 28688
rect 7009 28679 7067 28685
rect 7009 28645 7021 28679
rect 7055 28676 7067 28679
rect 10686 28676 10692 28688
rect 7055 28648 10692 28676
rect 7055 28645 7067 28648
rect 7009 28639 7067 28645
rect 10686 28636 10692 28648
rect 10744 28676 10750 28688
rect 12360 28676 12388 28707
rect 14550 28704 14556 28716
rect 14608 28704 14614 28756
rect 14642 28704 14648 28756
rect 14700 28744 14706 28756
rect 14737 28747 14795 28753
rect 14737 28744 14749 28747
rect 14700 28716 14749 28744
rect 14700 28704 14706 28716
rect 14737 28713 14749 28716
rect 14783 28713 14795 28747
rect 14737 28707 14795 28713
rect 19061 28747 19119 28753
rect 19061 28713 19073 28747
rect 19107 28744 19119 28747
rect 21177 28747 21235 28753
rect 19107 28716 20208 28744
rect 19107 28713 19119 28716
rect 19061 28707 19119 28713
rect 10744 28648 12388 28676
rect 14568 28676 14596 28704
rect 15105 28679 15163 28685
rect 15105 28676 15117 28679
rect 14568 28648 15117 28676
rect 10744 28636 10750 28648
rect 15105 28645 15117 28648
rect 15151 28645 15163 28679
rect 15105 28639 15163 28645
rect 19334 28636 19340 28688
rect 19392 28676 19398 28688
rect 20180 28685 20208 28716
rect 21177 28713 21189 28747
rect 21223 28744 21235 28747
rect 21450 28744 21456 28756
rect 21223 28716 21456 28744
rect 21223 28713 21235 28716
rect 21177 28707 21235 28713
rect 21450 28704 21456 28716
rect 21508 28704 21514 28756
rect 23474 28704 23480 28756
rect 23532 28744 23538 28756
rect 23661 28747 23719 28753
rect 23661 28744 23673 28747
rect 23532 28716 23673 28744
rect 23532 28704 23538 28716
rect 23661 28713 23673 28716
rect 23707 28713 23719 28747
rect 23661 28707 23719 28713
rect 25314 28704 25320 28756
rect 25372 28744 25378 28756
rect 25430 28747 25488 28753
rect 25430 28744 25442 28747
rect 25372 28716 25442 28744
rect 25372 28704 25378 28716
rect 25430 28713 25442 28716
rect 25476 28713 25488 28747
rect 25430 28707 25488 28713
rect 26099 28747 26157 28753
rect 26099 28713 26111 28747
rect 26145 28744 26157 28747
rect 26326 28744 26332 28756
rect 26145 28716 26332 28744
rect 26145 28713 26157 28716
rect 26099 28707 26157 28713
rect 26326 28704 26332 28716
rect 26384 28704 26390 28756
rect 28258 28704 28264 28756
rect 28316 28744 28322 28756
rect 28813 28747 28871 28753
rect 28813 28744 28825 28747
rect 28316 28716 28825 28744
rect 28316 28704 28322 28716
rect 28813 28713 28825 28716
rect 28859 28713 28871 28747
rect 28813 28707 28871 28713
rect 28994 28704 29000 28756
rect 29052 28744 29058 28756
rect 30653 28747 30711 28753
rect 30653 28744 30665 28747
rect 29052 28716 30665 28744
rect 29052 28704 29058 28716
rect 30653 28713 30665 28716
rect 30699 28713 30711 28747
rect 30653 28707 30711 28713
rect 19981 28679 20039 28685
rect 19981 28676 19993 28679
rect 19392 28648 19993 28676
rect 19392 28636 19398 28648
rect 19981 28645 19993 28648
rect 20027 28645 20039 28679
rect 19981 28639 20039 28645
rect 20165 28679 20223 28685
rect 20165 28645 20177 28679
rect 20211 28645 20223 28679
rect 22097 28679 22155 28685
rect 22097 28676 22109 28679
rect 20165 28639 20223 28645
rect 21284 28648 22109 28676
rect 1394 28568 1400 28620
rect 1452 28608 1458 28620
rect 1765 28611 1823 28617
rect 1765 28608 1777 28611
rect 1452 28580 1777 28608
rect 1452 28568 1458 28580
rect 1765 28577 1777 28580
rect 1811 28608 1823 28611
rect 3878 28608 3884 28620
rect 1811 28580 3884 28608
rect 1811 28577 1823 28580
rect 1765 28571 1823 28577
rect 3878 28568 3884 28580
rect 3936 28608 3942 28620
rect 4801 28611 4859 28617
rect 4801 28608 4813 28611
rect 3936 28580 4813 28608
rect 3936 28568 3942 28580
rect 4801 28577 4813 28580
rect 4847 28577 4859 28611
rect 4801 28571 4859 28577
rect 8294 28568 8300 28620
rect 8352 28608 8358 28620
rect 8389 28611 8447 28617
rect 8389 28608 8401 28611
rect 8352 28580 8401 28608
rect 8352 28568 8358 28580
rect 8389 28577 8401 28580
rect 8435 28577 8447 28611
rect 8570 28608 8576 28620
rect 8531 28580 8576 28608
rect 8389 28571 8447 28577
rect 5902 28500 5908 28552
rect 5960 28540 5966 28552
rect 7101 28543 7159 28549
rect 7101 28540 7113 28543
rect 5960 28512 7113 28540
rect 5960 28500 5966 28512
rect 7101 28509 7113 28512
rect 7147 28509 7159 28543
rect 7101 28503 7159 28509
rect 7285 28543 7343 28549
rect 7285 28509 7297 28543
rect 7331 28540 7343 28543
rect 7466 28540 7472 28552
rect 7331 28512 7472 28540
rect 7331 28509 7343 28512
rect 7285 28503 7343 28509
rect 7466 28500 7472 28512
rect 7524 28500 7530 28552
rect 8404 28540 8432 28571
rect 8570 28568 8576 28580
rect 8628 28568 8634 28620
rect 9674 28608 9680 28620
rect 9508 28580 9680 28608
rect 9508 28540 9536 28580
rect 9674 28568 9680 28580
rect 9732 28568 9738 28620
rect 9858 28608 9864 28620
rect 9819 28580 9864 28608
rect 9858 28568 9864 28580
rect 9916 28568 9922 28620
rect 10870 28568 10876 28620
rect 10928 28608 10934 28620
rect 10965 28611 11023 28617
rect 10965 28608 10977 28611
rect 10928 28580 10977 28608
rect 10928 28568 10934 28580
rect 10965 28577 10977 28580
rect 11011 28577 11023 28611
rect 10965 28571 11023 28577
rect 11054 28568 11060 28620
rect 11112 28608 11118 28620
rect 11221 28611 11279 28617
rect 11221 28608 11233 28611
rect 11112 28580 11233 28608
rect 11112 28568 11118 28580
rect 11221 28577 11233 28580
rect 11267 28577 11279 28611
rect 12802 28608 12808 28620
rect 12763 28580 12808 28608
rect 11221 28571 11279 28577
rect 12802 28568 12808 28580
rect 12860 28568 12866 28620
rect 12986 28608 12992 28620
rect 12947 28580 12992 28608
rect 12986 28568 12992 28580
rect 13044 28568 13050 28620
rect 13630 28608 13636 28620
rect 13543 28580 13636 28608
rect 13630 28568 13636 28580
rect 13688 28608 13694 28620
rect 13998 28608 14004 28620
rect 13688 28580 14004 28608
rect 13688 28568 13694 28580
rect 13998 28568 14004 28580
rect 14056 28568 14062 28620
rect 16758 28608 16764 28620
rect 16719 28580 16764 28608
rect 16758 28568 16764 28580
rect 16816 28568 16822 28620
rect 19058 28608 19064 28620
rect 19019 28580 19064 28608
rect 19058 28568 19064 28580
rect 19116 28568 19122 28620
rect 20254 28608 20260 28620
rect 20215 28580 20260 28608
rect 20254 28568 20260 28580
rect 20312 28568 20318 28620
rect 20901 28611 20959 28617
rect 20901 28577 20913 28611
rect 20947 28577 20959 28611
rect 20901 28571 20959 28577
rect 8404 28512 9536 28540
rect 9585 28543 9643 28549
rect 9585 28509 9597 28543
rect 9631 28540 9643 28543
rect 10042 28540 10048 28552
rect 9631 28512 10048 28540
rect 9631 28509 9643 28512
rect 9585 28503 9643 28509
rect 10042 28500 10048 28512
rect 10100 28500 10106 28552
rect 13725 28543 13783 28549
rect 13725 28509 13737 28543
rect 13771 28540 13783 28543
rect 15197 28543 15255 28549
rect 15197 28540 15209 28543
rect 13771 28512 15209 28540
rect 13771 28509 13783 28512
rect 13725 28503 13783 28509
rect 15197 28509 15209 28512
rect 15243 28509 15255 28543
rect 15197 28503 15255 28509
rect 15289 28543 15347 28549
rect 15289 28509 15301 28543
rect 15335 28509 15347 28543
rect 15289 28503 15347 28509
rect 16577 28543 16635 28549
rect 16577 28509 16589 28543
rect 16623 28540 16635 28543
rect 16666 28540 16672 28552
rect 16623 28512 16672 28540
rect 16623 28509 16635 28512
rect 16577 28503 16635 28509
rect 13354 28432 13360 28484
rect 13412 28472 13418 28484
rect 15304 28472 15332 28503
rect 16666 28500 16672 28512
rect 16724 28500 16730 28552
rect 18785 28543 18843 28549
rect 18785 28509 18797 28543
rect 18831 28540 18843 28543
rect 20346 28540 20352 28552
rect 18831 28512 20352 28540
rect 18831 28509 18843 28512
rect 18785 28503 18843 28509
rect 20346 28500 20352 28512
rect 20404 28500 20410 28552
rect 18966 28472 18972 28484
rect 13412 28444 15332 28472
rect 18927 28444 18972 28472
rect 13412 28432 13418 28444
rect 18966 28432 18972 28444
rect 19024 28432 19030 28484
rect 20916 28472 20944 28571
rect 20990 28568 20996 28620
rect 21048 28608 21054 28620
rect 21284 28617 21312 28648
rect 22097 28645 22109 28648
rect 22143 28645 22155 28679
rect 24762 28676 24768 28688
rect 22097 28639 22155 28645
rect 24044 28648 24768 28676
rect 21269 28611 21327 28617
rect 21048 28580 21093 28608
rect 21048 28568 21054 28580
rect 21269 28577 21281 28611
rect 21315 28577 21327 28611
rect 22002 28608 22008 28620
rect 21963 28580 22008 28608
rect 21269 28571 21327 28577
rect 22002 28568 22008 28580
rect 22060 28568 22066 28620
rect 22189 28611 22247 28617
rect 22189 28577 22201 28611
rect 22235 28608 22247 28611
rect 22554 28608 22560 28620
rect 22235 28580 22560 28608
rect 22235 28577 22247 28580
rect 22189 28571 22247 28577
rect 22554 28568 22560 28580
rect 22612 28568 22618 28620
rect 23937 28611 23995 28617
rect 23937 28577 23949 28611
rect 23983 28608 23995 28611
rect 24044 28608 24072 28648
rect 24762 28636 24768 28648
rect 24820 28676 24826 28688
rect 25225 28679 25283 28685
rect 25225 28676 25237 28679
rect 24820 28648 25237 28676
rect 24820 28636 24826 28648
rect 25225 28645 25237 28648
rect 25271 28645 25283 28679
rect 25225 28639 25283 28645
rect 26510 28636 26516 28688
rect 26568 28636 26574 28688
rect 29181 28679 29239 28685
rect 29181 28645 29193 28679
rect 29227 28676 29239 28679
rect 30282 28676 30288 28688
rect 29227 28648 30288 28676
rect 29227 28645 29239 28648
rect 29181 28639 29239 28645
rect 30282 28636 30288 28648
rect 30340 28636 30346 28688
rect 32398 28685 32404 28688
rect 32392 28676 32404 28685
rect 32359 28648 32404 28676
rect 32392 28639 32404 28648
rect 32398 28636 32404 28639
rect 32456 28636 32462 28688
rect 23983 28580 24072 28608
rect 24121 28611 24179 28617
rect 23983 28577 23995 28580
rect 23937 28571 23995 28577
rect 24121 28577 24133 28611
rect 24167 28608 24179 28611
rect 24302 28608 24308 28620
rect 24167 28580 24308 28608
rect 24167 28577 24179 28580
rect 24121 28571 24179 28577
rect 24302 28568 24308 28580
rect 24360 28568 24366 28620
rect 27614 28568 27620 28620
rect 27672 28608 27678 28620
rect 27893 28611 27951 28617
rect 27893 28608 27905 28611
rect 27672 28580 27905 28608
rect 27672 28568 27678 28580
rect 27893 28577 27905 28580
rect 27939 28577 27951 28611
rect 31021 28611 31079 28617
rect 31021 28608 31033 28611
rect 27893 28571 27951 28577
rect 29288 28580 31033 28608
rect 29288 28552 29316 28580
rect 31021 28577 31033 28580
rect 31067 28577 31079 28611
rect 31021 28571 31079 28577
rect 21082 28540 21088 28552
rect 21043 28512 21088 28540
rect 21082 28500 21088 28512
rect 21140 28500 21146 28552
rect 23845 28543 23903 28549
rect 23845 28509 23857 28543
rect 23891 28509 23903 28543
rect 23845 28503 23903 28509
rect 24029 28543 24087 28549
rect 24029 28509 24041 28543
rect 24075 28509 24087 28543
rect 24029 28503 24087 28509
rect 23860 28472 23888 28503
rect 23934 28472 23940 28484
rect 20916 28444 22876 28472
rect 23860 28444 23940 28472
rect 22848 28416 22876 28444
rect 23934 28432 23940 28444
rect 23992 28432 23998 28484
rect 6270 28364 6276 28416
rect 6328 28404 6334 28416
rect 6641 28407 6699 28413
rect 6641 28404 6653 28407
rect 6328 28376 6653 28404
rect 6328 28364 6334 28376
rect 6641 28373 6653 28376
rect 6687 28373 6699 28407
rect 6641 28367 6699 28373
rect 12618 28364 12624 28416
rect 12676 28404 12682 28416
rect 12897 28407 12955 28413
rect 12897 28404 12909 28407
rect 12676 28376 12909 28404
rect 12676 28364 12682 28376
rect 12897 28373 12909 28376
rect 12943 28373 12955 28407
rect 16942 28404 16948 28416
rect 16903 28376 16948 28404
rect 12897 28367 12955 28373
rect 16942 28364 16948 28376
rect 17000 28364 17006 28416
rect 19334 28364 19340 28416
rect 19392 28404 19398 28416
rect 20073 28407 20131 28413
rect 20073 28404 20085 28407
rect 19392 28376 20085 28404
rect 19392 28364 19398 28376
rect 20073 28373 20085 28376
rect 20119 28373 20131 28407
rect 20073 28367 20131 28373
rect 22830 28364 22836 28416
rect 22888 28404 22894 28416
rect 24044 28404 24072 28503
rect 25774 28500 25780 28552
rect 25832 28540 25838 28552
rect 27525 28543 27583 28549
rect 27525 28540 27537 28543
rect 25832 28512 27537 28540
rect 25832 28500 25838 28512
rect 27525 28509 27537 28512
rect 27571 28509 27583 28543
rect 29270 28540 29276 28552
rect 29231 28512 29276 28540
rect 27525 28503 27583 28509
rect 29270 28500 29276 28512
rect 29328 28500 29334 28552
rect 29457 28543 29515 28549
rect 29457 28509 29469 28543
rect 29503 28509 29515 28543
rect 29457 28503 29515 28509
rect 29472 28472 29500 28503
rect 30282 28500 30288 28552
rect 30340 28540 30346 28552
rect 30469 28543 30527 28549
rect 30469 28540 30481 28543
rect 30340 28512 30481 28540
rect 30340 28500 30346 28512
rect 30469 28509 30481 28512
rect 30515 28509 30527 28543
rect 30469 28503 30527 28509
rect 30929 28543 30987 28549
rect 30929 28509 30941 28543
rect 30975 28540 30987 28543
rect 31294 28540 31300 28552
rect 30975 28512 31300 28540
rect 30975 28509 30987 28512
rect 30929 28503 30987 28509
rect 31294 28500 31300 28512
rect 31352 28500 31358 28552
rect 31938 28500 31944 28552
rect 31996 28540 32002 28552
rect 32125 28543 32183 28549
rect 32125 28540 32137 28543
rect 31996 28512 32137 28540
rect 31996 28500 32002 28512
rect 32125 28509 32137 28512
rect 32171 28509 32183 28543
rect 32125 28503 32183 28509
rect 31202 28472 31208 28484
rect 29472 28444 31208 28472
rect 31202 28432 31208 28444
rect 31260 28432 31266 28484
rect 22888 28376 24072 28404
rect 22888 28364 22894 28376
rect 24118 28364 24124 28416
rect 24176 28404 24182 28416
rect 25222 28404 25228 28416
rect 24176 28376 25228 28404
rect 24176 28364 24182 28376
rect 25222 28364 25228 28376
rect 25280 28404 25286 28416
rect 25409 28407 25467 28413
rect 25409 28404 25421 28407
rect 25280 28376 25421 28404
rect 25280 28364 25286 28376
rect 25409 28373 25421 28376
rect 25455 28373 25467 28407
rect 25409 28367 25467 28373
rect 25593 28407 25651 28413
rect 25593 28373 25605 28407
rect 25639 28404 25651 28407
rect 25682 28404 25688 28416
rect 25639 28376 25688 28404
rect 25639 28373 25651 28376
rect 25593 28367 25651 28373
rect 25682 28364 25688 28376
rect 25740 28364 25746 28416
rect 33502 28404 33508 28416
rect 33463 28376 33508 28404
rect 33502 28364 33508 28376
rect 33560 28364 33566 28416
rect 1104 28314 34316 28336
rect 1104 28262 6517 28314
rect 6569 28262 6581 28314
rect 6633 28262 6645 28314
rect 6697 28262 6709 28314
rect 6761 28262 17588 28314
rect 17640 28262 17652 28314
rect 17704 28262 17716 28314
rect 17768 28262 17780 28314
rect 17832 28262 28658 28314
rect 28710 28262 28722 28314
rect 28774 28262 28786 28314
rect 28838 28262 28850 28314
rect 28902 28262 34316 28314
rect 1104 28240 34316 28262
rect 3326 28160 3332 28212
rect 3384 28200 3390 28212
rect 3697 28203 3755 28209
rect 3697 28200 3709 28203
rect 3384 28172 3709 28200
rect 3384 28160 3390 28172
rect 3697 28169 3709 28172
rect 3743 28169 3755 28203
rect 4430 28200 4436 28212
rect 4391 28172 4436 28200
rect 3697 28163 3755 28169
rect 4430 28160 4436 28172
rect 4488 28160 4494 28212
rect 5534 28200 5540 28212
rect 5495 28172 5540 28200
rect 5534 28160 5540 28172
rect 5592 28160 5598 28212
rect 11054 28200 11060 28212
rect 11015 28172 11060 28200
rect 11054 28160 11060 28172
rect 11112 28160 11118 28212
rect 12989 28203 13047 28209
rect 12989 28169 13001 28203
rect 13035 28200 13047 28203
rect 13906 28200 13912 28212
rect 13035 28172 13912 28200
rect 13035 28169 13047 28172
rect 12989 28163 13047 28169
rect 13906 28160 13912 28172
rect 13964 28160 13970 28212
rect 20257 28203 20315 28209
rect 20257 28169 20269 28203
rect 20303 28200 20315 28203
rect 21082 28200 21088 28212
rect 20303 28172 21088 28200
rect 20303 28169 20315 28172
rect 20257 28163 20315 28169
rect 21082 28160 21088 28172
rect 21140 28160 21146 28212
rect 25774 28200 25780 28212
rect 25735 28172 25780 28200
rect 25774 28160 25780 28172
rect 25832 28160 25838 28212
rect 29270 28160 29276 28212
rect 29328 28200 29334 28212
rect 30193 28203 30251 28209
rect 30193 28200 30205 28203
rect 29328 28172 30205 28200
rect 29328 28160 29334 28172
rect 30193 28169 30205 28172
rect 30239 28169 30251 28203
rect 30193 28163 30251 28169
rect 17310 28092 17316 28144
rect 17368 28132 17374 28144
rect 17405 28135 17463 28141
rect 17405 28132 17417 28135
rect 17368 28104 17417 28132
rect 17368 28092 17374 28104
rect 17405 28101 17417 28104
rect 17451 28101 17463 28135
rect 20901 28135 20959 28141
rect 20901 28132 20913 28135
rect 17405 28095 17463 28101
rect 20180 28104 20913 28132
rect 9490 28024 9496 28076
rect 9548 28064 9554 28076
rect 9861 28067 9919 28073
rect 9861 28064 9873 28067
rect 9548 28036 9873 28064
rect 9548 28024 9554 28036
rect 9861 28033 9873 28036
rect 9907 28033 9919 28067
rect 9861 28027 9919 28033
rect 13722 28024 13728 28076
rect 13780 28064 13786 28076
rect 14737 28067 14795 28073
rect 14737 28064 14749 28067
rect 13780 28036 14749 28064
rect 13780 28024 13786 28036
rect 14737 28033 14749 28036
rect 14783 28033 14795 28067
rect 14737 28027 14795 28033
rect 16942 28024 16948 28076
rect 17000 28064 17006 28076
rect 17773 28067 17831 28073
rect 17773 28064 17785 28067
rect 17000 28036 17785 28064
rect 17000 28024 17006 28036
rect 17773 28033 17785 28036
rect 17819 28033 17831 28067
rect 19150 28064 19156 28076
rect 19111 28036 19156 28064
rect 17773 28027 17831 28033
rect 19150 28024 19156 28036
rect 19208 28024 19214 28076
rect 20180 28064 20208 28104
rect 20901 28101 20913 28104
rect 20947 28101 20959 28135
rect 20901 28095 20959 28101
rect 24949 28135 25007 28141
rect 24949 28101 24961 28135
rect 24995 28132 25007 28135
rect 25547 28135 25605 28141
rect 25547 28132 25559 28135
rect 24995 28104 25559 28132
rect 24995 28101 25007 28104
rect 24949 28095 25007 28101
rect 25547 28101 25559 28104
rect 25593 28101 25605 28135
rect 25682 28132 25688 28144
rect 25643 28104 25688 28132
rect 25547 28095 25605 28101
rect 25682 28092 25688 28104
rect 25740 28092 25746 28144
rect 20254 28064 20260 28076
rect 20180 28036 20260 28064
rect 5353 27999 5411 28005
rect 5353 27965 5365 27999
rect 5399 27996 5411 27999
rect 6270 27996 6276 28008
rect 5399 27968 6276 27996
rect 5399 27965 5411 27968
rect 5353 27959 5411 27965
rect 6270 27956 6276 27968
rect 6328 27956 6334 28008
rect 8113 27999 8171 28005
rect 8113 27965 8125 27999
rect 8159 27996 8171 27999
rect 8202 27996 8208 28008
rect 8159 27968 8208 27996
rect 8159 27965 8171 27968
rect 8113 27959 8171 27965
rect 8202 27956 8208 27968
rect 8260 27956 8266 28008
rect 8297 27999 8355 28005
rect 8297 27965 8309 27999
rect 8343 27996 8355 27999
rect 8386 27996 8392 28008
rect 8343 27968 8392 27996
rect 8343 27965 8355 27968
rect 8297 27959 8355 27965
rect 8386 27956 8392 27968
rect 8444 27956 8450 28008
rect 10045 27999 10103 28005
rect 10045 27965 10057 27999
rect 10091 27965 10103 27999
rect 10226 27996 10232 28008
rect 10187 27968 10232 27996
rect 10045 27959 10103 27965
rect 2958 27888 2964 27940
rect 3016 27928 3022 27940
rect 3605 27931 3663 27937
rect 3605 27928 3617 27931
rect 3016 27900 3617 27928
rect 3016 27888 3022 27900
rect 3605 27897 3617 27900
rect 3651 27897 3663 27931
rect 4338 27928 4344 27940
rect 4299 27900 4344 27928
rect 3605 27891 3663 27897
rect 4338 27888 4344 27900
rect 4396 27928 4402 27940
rect 5169 27931 5227 27937
rect 5169 27928 5181 27931
rect 4396 27900 5181 27928
rect 4396 27888 4402 27900
rect 5169 27897 5181 27900
rect 5215 27897 5227 27931
rect 10060 27928 10088 27959
rect 10226 27956 10232 27968
rect 10284 27956 10290 28008
rect 10962 27996 10968 28008
rect 10923 27968 10968 27996
rect 10962 27956 10968 27968
rect 11020 27956 11026 28008
rect 11149 27999 11207 28005
rect 11149 27965 11161 27999
rect 11195 27996 11207 27999
rect 12618 27996 12624 28008
rect 11195 27968 12624 27996
rect 11195 27965 11207 27968
rect 11149 27959 11207 27965
rect 12618 27956 12624 27968
rect 12676 27956 12682 28008
rect 12805 27999 12863 28005
rect 12805 27965 12817 27999
rect 12851 27965 12863 27999
rect 12805 27959 12863 27965
rect 12989 27999 13047 28005
rect 12989 27965 13001 27999
rect 13035 27996 13047 27999
rect 13078 27996 13084 28008
rect 13035 27968 13084 27996
rect 13035 27965 13047 27968
rect 12989 27959 13047 27965
rect 10134 27928 10140 27940
rect 10060 27900 10140 27928
rect 5169 27891 5227 27897
rect 10134 27888 10140 27900
rect 10192 27888 10198 27940
rect 12342 27888 12348 27940
rect 12400 27928 12406 27940
rect 12820 27928 12848 27959
rect 13078 27956 13084 27968
rect 13136 27956 13142 28008
rect 14645 27999 14703 28005
rect 14645 27965 14657 27999
rect 14691 27996 14703 27999
rect 15010 27996 15016 28008
rect 14691 27968 15016 27996
rect 14691 27965 14703 27968
rect 14645 27959 14703 27965
rect 15010 27956 15016 27968
rect 15068 27956 15074 28008
rect 20180 28005 20208 28036
rect 20254 28024 20260 28036
rect 20312 28024 20318 28076
rect 20438 28064 20444 28076
rect 20351 28036 20444 28064
rect 20364 28005 20392 28036
rect 20438 28024 20444 28036
rect 20496 28064 20502 28076
rect 21545 28067 21603 28073
rect 21545 28064 21557 28067
rect 20496 28036 21557 28064
rect 20496 28024 20502 28036
rect 21545 28033 21557 28036
rect 21591 28033 21603 28067
rect 24854 28064 24860 28076
rect 21545 28027 21603 28033
rect 23952 28036 24860 28064
rect 18877 27999 18935 28005
rect 18877 27965 18889 27999
rect 18923 27996 18935 27999
rect 20165 27999 20223 28005
rect 20165 27996 20177 27999
rect 18923 27968 20177 27996
rect 18923 27965 18935 27968
rect 18877 27959 18935 27965
rect 20165 27965 20177 27968
rect 20211 27965 20223 27999
rect 20165 27959 20223 27965
rect 20349 27999 20407 28005
rect 20349 27965 20361 27999
rect 20395 27965 20407 27999
rect 20806 27996 20812 28008
rect 20767 27968 20812 27996
rect 20349 27959 20407 27965
rect 20806 27956 20812 27968
rect 20864 27956 20870 28008
rect 20993 27999 21051 28005
rect 20993 27965 21005 27999
rect 21039 27996 21051 27999
rect 21082 27996 21088 28008
rect 21039 27968 21088 27996
rect 21039 27965 21051 27968
rect 20993 27959 21051 27965
rect 21082 27956 21088 27968
rect 21140 27956 21146 28008
rect 23952 28005 23980 28036
rect 24854 28024 24860 28036
rect 24912 28024 24918 28076
rect 26421 28067 26479 28073
rect 26421 28064 26433 28067
rect 25884 28036 26433 28064
rect 21453 27999 21511 28005
rect 21453 27965 21465 27999
rect 21499 27965 21511 27999
rect 23937 27999 23995 28005
rect 21453 27959 21511 27965
rect 22066 27968 23888 27996
rect 17954 27928 17960 27940
rect 12400 27900 12848 27928
rect 17915 27900 17960 27928
rect 12400 27888 12406 27900
rect 17954 27888 17960 27900
rect 18012 27888 18018 27940
rect 20714 27888 20720 27940
rect 20772 27928 20778 27940
rect 21468 27928 21496 27959
rect 20772 27900 21496 27928
rect 20772 27888 20778 27900
rect 8202 27860 8208 27872
rect 8163 27832 8208 27860
rect 8202 27820 8208 27832
rect 8260 27820 8266 27872
rect 14182 27860 14188 27872
rect 14143 27832 14188 27860
rect 14182 27820 14188 27832
rect 14240 27820 14246 27872
rect 14550 27860 14556 27872
rect 14511 27832 14556 27860
rect 14550 27820 14556 27832
rect 14608 27820 14614 27872
rect 17402 27820 17408 27872
rect 17460 27860 17466 27872
rect 17865 27863 17923 27869
rect 17865 27860 17877 27863
rect 17460 27832 17877 27860
rect 17460 27820 17466 27832
rect 17865 27829 17877 27832
rect 17911 27829 17923 27863
rect 18506 27860 18512 27872
rect 18467 27832 18512 27860
rect 17865 27823 17923 27829
rect 18506 27820 18512 27832
rect 18564 27820 18570 27872
rect 18969 27863 19027 27869
rect 18969 27829 18981 27863
rect 19015 27860 19027 27863
rect 19058 27860 19064 27872
rect 19015 27832 19064 27860
rect 19015 27829 19027 27832
rect 18969 27823 19027 27829
rect 19058 27820 19064 27832
rect 19116 27820 19122 27872
rect 19150 27820 19156 27872
rect 19208 27860 19214 27872
rect 21174 27860 21180 27872
rect 19208 27832 21180 27860
rect 19208 27820 19214 27832
rect 21174 27820 21180 27832
rect 21232 27860 21238 27872
rect 22066 27860 22094 27968
rect 22554 27888 22560 27940
rect 22612 27928 22618 27940
rect 23017 27931 23075 27937
rect 23017 27928 23029 27931
rect 22612 27900 23029 27928
rect 22612 27888 22618 27900
rect 23017 27897 23029 27900
rect 23063 27897 23075 27931
rect 23017 27891 23075 27897
rect 21232 27832 22094 27860
rect 21232 27820 21238 27832
rect 22830 27820 22836 27872
rect 22888 27860 22894 27872
rect 23109 27863 23167 27869
rect 23109 27860 23121 27863
rect 22888 27832 23121 27860
rect 22888 27820 22894 27832
rect 23109 27829 23121 27832
rect 23155 27829 23167 27863
rect 23109 27823 23167 27829
rect 23566 27820 23572 27872
rect 23624 27860 23630 27872
rect 23753 27863 23811 27869
rect 23753 27860 23765 27863
rect 23624 27832 23765 27860
rect 23624 27820 23630 27832
rect 23753 27829 23765 27832
rect 23799 27829 23811 27863
rect 23860 27860 23888 27968
rect 23937 27965 23949 27999
rect 23983 27965 23995 27999
rect 23937 27959 23995 27965
rect 24026 27956 24032 28008
rect 24084 27996 24090 28008
rect 24213 27999 24271 28005
rect 24213 27996 24225 27999
rect 24084 27968 24225 27996
rect 24084 27956 24090 27968
rect 24213 27965 24225 27968
rect 24259 27996 24271 27999
rect 24673 27999 24731 28005
rect 24673 27996 24685 27999
rect 24259 27968 24685 27996
rect 24259 27965 24271 27968
rect 24213 27959 24271 27965
rect 24673 27965 24685 27968
rect 24719 27965 24731 27999
rect 24673 27959 24731 27965
rect 24762 27956 24768 28008
rect 24820 27996 24826 28008
rect 24949 27999 25007 28005
rect 24820 27968 24865 27996
rect 24820 27956 24826 27968
rect 24949 27965 24961 27999
rect 24995 27996 25007 27999
rect 25314 27996 25320 28008
rect 24995 27968 25320 27996
rect 24995 27965 25007 27968
rect 24949 27959 25007 27965
rect 25314 27956 25320 27968
rect 25372 27956 25378 28008
rect 25884 28005 25912 28036
rect 26421 28033 26433 28036
rect 26467 28033 26479 28067
rect 26421 28027 26479 28033
rect 27614 28024 27620 28076
rect 27672 28064 27678 28076
rect 28445 28067 28503 28073
rect 28445 28064 28457 28067
rect 27672 28036 28457 28064
rect 27672 28024 27678 28036
rect 28445 28033 28457 28036
rect 28491 28033 28503 28067
rect 28445 28027 28503 28033
rect 25409 27999 25467 28005
rect 25409 27965 25421 27999
rect 25455 27965 25467 27999
rect 25409 27959 25467 27965
rect 25869 27999 25927 28005
rect 25869 27965 25881 27999
rect 25915 27965 25927 27999
rect 26326 27996 26332 28008
rect 26287 27968 26332 27996
rect 25869 27959 25927 27965
rect 24121 27931 24179 27937
rect 24121 27897 24133 27931
rect 24167 27928 24179 27931
rect 24780 27928 24808 27956
rect 24167 27900 24808 27928
rect 25424 27928 25452 27959
rect 26326 27956 26332 27968
rect 26384 27956 26390 28008
rect 26513 27999 26571 28005
rect 26513 27965 26525 27999
rect 26559 27996 26571 27999
rect 26602 27996 26608 28008
rect 26559 27968 26608 27996
rect 26559 27965 26571 27968
rect 26513 27959 26571 27965
rect 26602 27956 26608 27968
rect 26660 27956 26666 28008
rect 30208 27996 30236 28163
rect 31202 28160 31208 28212
rect 31260 28200 31266 28212
rect 31665 28203 31723 28209
rect 31665 28200 31677 28203
rect 31260 28172 31677 28200
rect 31260 28160 31266 28172
rect 31665 28169 31677 28172
rect 31711 28169 31723 28203
rect 31665 28163 31723 28169
rect 30837 27999 30895 28005
rect 30837 27996 30849 27999
rect 30208 27968 30849 27996
rect 30837 27965 30849 27968
rect 30883 27965 30895 27999
rect 30837 27959 30895 27965
rect 31021 27999 31079 28005
rect 31021 27965 31033 27999
rect 31067 27996 31079 27999
rect 31481 27999 31539 28005
rect 31481 27996 31493 27999
rect 31067 27968 31493 27996
rect 31067 27965 31079 27968
rect 31021 27959 31079 27965
rect 31481 27965 31493 27968
rect 31527 27965 31539 27999
rect 31481 27959 31539 27965
rect 26050 27928 26056 27940
rect 25424 27900 26056 27928
rect 24167 27897 24179 27900
rect 24121 27891 24179 27897
rect 26050 27888 26056 27900
rect 26108 27888 26114 27940
rect 28718 27928 28724 27940
rect 28679 27900 28724 27928
rect 28718 27888 28724 27900
rect 28776 27888 28782 27940
rect 30098 27928 30104 27940
rect 29946 27900 30104 27928
rect 30098 27888 30104 27900
rect 30156 27888 30162 27940
rect 30374 27888 30380 27940
rect 30432 27928 30438 27940
rect 31036 27928 31064 27959
rect 30432 27900 31064 27928
rect 30432 27888 30438 27900
rect 25774 27860 25780 27872
rect 23860 27832 25780 27860
rect 23753 27823 23811 27829
rect 25774 27820 25780 27832
rect 25832 27820 25838 27872
rect 30650 27860 30656 27872
rect 30611 27832 30656 27860
rect 30650 27820 30656 27832
rect 30708 27820 30714 27872
rect 1104 27770 34316 27792
rect 1104 27718 12052 27770
rect 12104 27718 12116 27770
rect 12168 27718 12180 27770
rect 12232 27718 12244 27770
rect 12296 27718 23123 27770
rect 23175 27718 23187 27770
rect 23239 27718 23251 27770
rect 23303 27718 23315 27770
rect 23367 27718 34316 27770
rect 1104 27696 34316 27718
rect 4246 27616 4252 27668
rect 4304 27656 4310 27668
rect 4709 27659 4767 27665
rect 4709 27656 4721 27659
rect 4304 27628 4721 27656
rect 4304 27616 4310 27628
rect 4709 27625 4721 27628
rect 4755 27625 4767 27659
rect 4709 27619 4767 27625
rect 12986 27616 12992 27668
rect 13044 27656 13050 27668
rect 13081 27659 13139 27665
rect 13081 27656 13093 27659
rect 13044 27628 13093 27656
rect 13044 27616 13050 27628
rect 13081 27625 13093 27628
rect 13127 27625 13139 27659
rect 13081 27619 13139 27625
rect 14550 27616 14556 27668
rect 14608 27656 14614 27668
rect 14737 27659 14795 27665
rect 14737 27656 14749 27659
rect 14608 27628 14749 27656
rect 14608 27616 14614 27628
rect 14737 27625 14749 27628
rect 14783 27625 14795 27659
rect 14737 27619 14795 27625
rect 15010 27616 15016 27668
rect 15068 27656 15074 27668
rect 15105 27659 15163 27665
rect 15105 27656 15117 27659
rect 15068 27628 15117 27656
rect 15068 27616 15074 27628
rect 15105 27625 15117 27628
rect 15151 27625 15163 27659
rect 20990 27656 20996 27668
rect 20951 27628 20996 27656
rect 15105 27619 15163 27625
rect 20990 27616 20996 27628
rect 21048 27616 21054 27668
rect 22094 27656 22100 27668
rect 21652 27628 22100 27656
rect 10045 27591 10103 27597
rect 10045 27557 10057 27591
rect 10091 27588 10103 27591
rect 10134 27588 10140 27600
rect 10091 27560 10140 27588
rect 10091 27557 10103 27560
rect 10045 27551 10103 27557
rect 10134 27548 10140 27560
rect 10192 27548 10198 27600
rect 10410 27588 10416 27600
rect 10371 27560 10416 27588
rect 10410 27548 10416 27560
rect 10468 27548 10474 27600
rect 11422 27588 11428 27600
rect 11383 27560 11428 27588
rect 11422 27548 11428 27560
rect 11480 27548 11486 27600
rect 13541 27591 13599 27597
rect 13541 27557 13553 27591
rect 13587 27588 13599 27591
rect 14182 27588 14188 27600
rect 13587 27560 14188 27588
rect 13587 27557 13599 27560
rect 13541 27551 13599 27557
rect 14182 27548 14188 27560
rect 14240 27548 14246 27600
rect 18414 27548 18420 27600
rect 18472 27548 18478 27600
rect 20714 27588 20720 27600
rect 20675 27560 20720 27588
rect 20714 27548 20720 27560
rect 20772 27548 20778 27600
rect 21652 27597 21680 27628
rect 22094 27616 22100 27628
rect 22152 27616 22158 27668
rect 25222 27656 25228 27668
rect 25183 27628 25228 27656
rect 25222 27616 25228 27628
rect 25280 27616 25286 27668
rect 28718 27616 28724 27668
rect 28776 27656 28782 27668
rect 28813 27659 28871 27665
rect 28813 27656 28825 27659
rect 28776 27628 28825 27656
rect 28776 27616 28782 27628
rect 28813 27625 28825 27628
rect 28859 27625 28871 27659
rect 32564 27659 32622 27665
rect 32564 27656 32576 27659
rect 28813 27619 28871 27625
rect 31726 27628 32576 27656
rect 31726 27597 31754 27628
rect 32564 27625 32576 27628
rect 32610 27656 32622 27659
rect 33502 27656 33508 27668
rect 32610 27628 33508 27656
rect 32610 27625 32622 27628
rect 32564 27619 32622 27625
rect 33502 27616 33508 27628
rect 33560 27616 33566 27668
rect 21637 27591 21695 27597
rect 21637 27557 21649 27591
rect 21683 27557 21695 27591
rect 31696 27591 31754 27597
rect 21637 27551 21695 27557
rect 21744 27560 22508 27588
rect 2958 27520 2964 27532
rect 2919 27492 2964 27520
rect 2958 27480 2964 27492
rect 3016 27480 3022 27532
rect 4617 27523 4675 27529
rect 4617 27489 4629 27523
rect 4663 27489 4675 27523
rect 4617 27483 4675 27489
rect 7213 27523 7271 27529
rect 7213 27489 7225 27523
rect 7259 27520 7271 27523
rect 8205 27523 8263 27529
rect 7259 27492 7604 27520
rect 7259 27489 7271 27492
rect 7213 27483 7271 27489
rect 2774 27412 2780 27464
rect 2832 27452 2838 27464
rect 2869 27455 2927 27461
rect 2869 27452 2881 27455
rect 2832 27424 2881 27452
rect 2832 27412 2838 27424
rect 2869 27421 2881 27424
rect 2915 27421 2927 27455
rect 2869 27415 2927 27421
rect 3053 27455 3111 27461
rect 3053 27421 3065 27455
rect 3099 27421 3111 27455
rect 3053 27415 3111 27421
rect 3068 27384 3096 27415
rect 3142 27412 3148 27464
rect 3200 27452 3206 27464
rect 3200 27424 3245 27452
rect 3200 27412 3206 27424
rect 4249 27387 4307 27393
rect 4249 27384 4261 27387
rect 3068 27356 4261 27384
rect 4249 27353 4261 27356
rect 4295 27353 4307 27387
rect 4632 27384 4660 27483
rect 4893 27455 4951 27461
rect 4893 27421 4905 27455
rect 4939 27452 4951 27455
rect 4982 27452 4988 27464
rect 4939 27424 4988 27452
rect 4939 27421 4951 27424
rect 4893 27415 4951 27421
rect 4982 27412 4988 27424
rect 5040 27412 5046 27464
rect 7469 27455 7527 27461
rect 7469 27421 7481 27455
rect 7515 27421 7527 27455
rect 7469 27415 7527 27421
rect 6086 27384 6092 27396
rect 4632 27356 6092 27384
rect 4249 27347 4307 27353
rect 6086 27344 6092 27356
rect 6144 27344 6150 27396
rect 2682 27316 2688 27328
rect 2643 27288 2688 27316
rect 2682 27276 2688 27288
rect 2740 27276 2746 27328
rect 4522 27276 4528 27328
rect 4580 27316 4586 27328
rect 7282 27316 7288 27328
rect 4580 27288 7288 27316
rect 4580 27276 4586 27288
rect 7282 27276 7288 27288
rect 7340 27316 7346 27328
rect 7484 27316 7512 27415
rect 7576 27384 7604 27492
rect 8205 27489 8217 27523
rect 8251 27489 8263 27523
rect 8386 27520 8392 27532
rect 8347 27492 8392 27520
rect 8205 27483 8263 27489
rect 8220 27452 8248 27483
rect 8386 27480 8392 27492
rect 8444 27480 8450 27532
rect 8481 27523 8539 27529
rect 8481 27489 8493 27523
rect 8527 27520 8539 27523
rect 9950 27520 9956 27532
rect 8527 27492 9956 27520
rect 8527 27489 8539 27492
rect 8481 27483 8539 27489
rect 9950 27480 9956 27492
rect 10008 27480 10014 27532
rect 10226 27520 10232 27532
rect 10187 27492 10232 27520
rect 10226 27480 10232 27492
rect 10284 27480 10290 27532
rect 11238 27480 11244 27532
rect 11296 27520 11302 27532
rect 11333 27523 11391 27529
rect 11333 27520 11345 27523
rect 11296 27492 11345 27520
rect 11296 27480 11302 27492
rect 11333 27489 11345 27492
rect 11379 27489 11391 27523
rect 11514 27520 11520 27532
rect 11475 27492 11520 27520
rect 11333 27483 11391 27489
rect 11514 27480 11520 27492
rect 11572 27480 11578 27532
rect 11698 27480 11704 27532
rect 11756 27520 11762 27532
rect 11977 27523 12035 27529
rect 11977 27520 11989 27523
rect 11756 27492 11989 27520
rect 11756 27480 11762 27492
rect 11977 27489 11989 27492
rect 12023 27489 12035 27523
rect 11977 27483 12035 27489
rect 12161 27523 12219 27529
rect 12161 27489 12173 27523
rect 12207 27520 12219 27523
rect 12434 27520 12440 27532
rect 12207 27492 12440 27520
rect 12207 27489 12219 27492
rect 12161 27483 12219 27489
rect 12434 27480 12440 27492
rect 12492 27480 12498 27532
rect 13446 27520 13452 27532
rect 13407 27492 13452 27520
rect 13446 27480 13452 27492
rect 13504 27480 13510 27532
rect 15010 27480 15016 27532
rect 15068 27520 15074 27532
rect 17218 27520 17224 27532
rect 15068 27492 15332 27520
rect 17179 27492 17224 27520
rect 15068 27480 15074 27492
rect 8754 27452 8760 27464
rect 8220 27424 8760 27452
rect 8754 27412 8760 27424
rect 8812 27412 8818 27464
rect 10042 27412 10048 27464
rect 10100 27452 10106 27464
rect 11054 27452 11060 27464
rect 10100 27424 11060 27452
rect 10100 27412 10106 27424
rect 11054 27412 11060 27424
rect 11112 27452 11118 27464
rect 11606 27452 11612 27464
rect 11112 27424 11612 27452
rect 11112 27412 11118 27424
rect 11606 27412 11612 27424
rect 11664 27452 11670 27464
rect 13633 27455 13691 27461
rect 13633 27452 13645 27455
rect 11664 27424 13645 27452
rect 11664 27412 11670 27424
rect 13633 27421 13645 27424
rect 13679 27452 13691 27455
rect 14734 27452 14740 27464
rect 13679 27424 14740 27452
rect 13679 27421 13691 27424
rect 13633 27415 13691 27421
rect 14734 27412 14740 27424
rect 14792 27412 14798 27464
rect 15304 27461 15332 27492
rect 17218 27480 17224 27492
rect 17276 27480 17282 27532
rect 18432 27520 18460 27548
rect 19426 27520 19432 27532
rect 18432 27492 19432 27520
rect 19426 27480 19432 27492
rect 19484 27480 19490 27532
rect 19794 27480 19800 27532
rect 19852 27520 19858 27532
rect 19981 27523 20039 27529
rect 19981 27520 19993 27523
rect 19852 27492 19993 27520
rect 19852 27480 19858 27492
rect 19981 27489 19993 27492
rect 20027 27489 20039 27523
rect 19981 27483 20039 27489
rect 20806 27480 20812 27532
rect 20864 27520 20870 27532
rect 20901 27523 20959 27529
rect 20901 27520 20913 27523
rect 20864 27492 20913 27520
rect 20864 27480 20870 27492
rect 20901 27489 20913 27492
rect 20947 27489 20959 27523
rect 20901 27483 20959 27489
rect 20993 27523 21051 27529
rect 20993 27489 21005 27523
rect 21039 27520 21051 27523
rect 21082 27520 21088 27532
rect 21039 27492 21088 27520
rect 21039 27489 21051 27492
rect 20993 27483 21051 27489
rect 15197 27455 15255 27461
rect 15197 27452 15209 27455
rect 15120 27424 15209 27452
rect 15120 27396 15148 27424
rect 15197 27421 15209 27424
rect 15243 27421 15255 27455
rect 15197 27415 15255 27421
rect 15289 27455 15347 27461
rect 15289 27421 15301 27455
rect 15335 27421 15347 27455
rect 15289 27415 15347 27421
rect 17589 27455 17647 27461
rect 17589 27421 17601 27455
rect 17635 27452 17647 27455
rect 18506 27452 18512 27464
rect 17635 27424 18512 27452
rect 17635 27421 17647 27424
rect 17589 27415 17647 27421
rect 18506 27412 18512 27424
rect 18564 27412 18570 27464
rect 20916 27452 20944 27483
rect 21082 27480 21088 27492
rect 21140 27520 21146 27532
rect 21744 27520 21772 27560
rect 21928 27529 21956 27560
rect 22480 27532 22508 27560
rect 31696 27557 31708 27591
rect 31742 27557 31754 27591
rect 31696 27551 31754 27557
rect 32769 27591 32827 27597
rect 32769 27557 32781 27591
rect 32815 27588 32827 27591
rect 33318 27588 33324 27600
rect 32815 27560 33324 27588
rect 32815 27557 32827 27560
rect 32769 27551 32827 27557
rect 33318 27548 33324 27560
rect 33376 27548 33382 27600
rect 21140 27492 21772 27520
rect 21821 27523 21879 27529
rect 21140 27480 21146 27492
rect 21821 27489 21833 27523
rect 21867 27489 21879 27523
rect 21821 27483 21879 27489
rect 21911 27523 21969 27529
rect 21911 27489 21923 27523
rect 21957 27489 21969 27523
rect 22370 27520 22376 27532
rect 21911 27483 21969 27489
rect 22020 27492 22376 27520
rect 21836 27452 21864 27483
rect 22020 27452 22048 27492
rect 22370 27480 22376 27492
rect 22428 27480 22434 27532
rect 22462 27480 22468 27532
rect 22520 27520 22526 27532
rect 22649 27523 22707 27529
rect 22520 27492 22565 27520
rect 22520 27480 22526 27492
rect 22649 27489 22661 27523
rect 22695 27489 22707 27523
rect 22649 27483 22707 27489
rect 24397 27523 24455 27529
rect 24397 27489 24409 27523
rect 24443 27520 24455 27523
rect 25038 27520 25044 27532
rect 24443 27492 25044 27520
rect 24443 27489 24455 27492
rect 24397 27483 24455 27489
rect 20916 27424 22048 27452
rect 22094 27412 22100 27464
rect 22152 27452 22158 27464
rect 22664 27452 22692 27483
rect 25038 27480 25044 27492
rect 25096 27480 25102 27532
rect 25130 27480 25136 27532
rect 25188 27520 25194 27532
rect 25225 27523 25283 27529
rect 25225 27520 25237 27523
rect 25188 27492 25237 27520
rect 25188 27480 25194 27492
rect 25225 27489 25237 27492
rect 25271 27489 25283 27523
rect 25225 27483 25283 27489
rect 25409 27523 25467 27529
rect 25409 27489 25421 27523
rect 25455 27520 25467 27523
rect 26234 27520 26240 27532
rect 25455 27492 26240 27520
rect 25455 27489 25467 27492
rect 25409 27483 25467 27489
rect 26234 27480 26240 27492
rect 26292 27520 26298 27532
rect 26694 27520 26700 27532
rect 26292 27492 26700 27520
rect 26292 27480 26298 27492
rect 26694 27480 26700 27492
rect 26752 27480 26758 27532
rect 28258 27480 28264 27532
rect 28316 27520 28322 27532
rect 28997 27523 29055 27529
rect 28997 27520 29009 27523
rect 28316 27492 29009 27520
rect 28316 27480 28322 27492
rect 28997 27489 29009 27492
rect 29043 27489 29055 27523
rect 28997 27483 29055 27489
rect 29273 27523 29331 27529
rect 29273 27489 29285 27523
rect 29319 27520 29331 27523
rect 30650 27520 30656 27532
rect 29319 27492 30656 27520
rect 29319 27489 29331 27492
rect 29273 27483 29331 27489
rect 30650 27480 30656 27492
rect 30708 27480 30714 27532
rect 31938 27452 31944 27464
rect 22152 27424 22692 27452
rect 31899 27424 31944 27452
rect 22152 27412 22158 27424
rect 31938 27412 31944 27424
rect 31996 27412 32002 27464
rect 8205 27387 8263 27393
rect 8205 27384 8217 27387
rect 7576 27356 8217 27384
rect 8205 27353 8217 27356
rect 8251 27353 8263 27387
rect 8205 27347 8263 27353
rect 15102 27344 15108 27396
rect 15160 27344 15166 27396
rect 24026 27384 24032 27396
rect 20180 27356 24032 27384
rect 20180 27328 20208 27356
rect 24026 27344 24032 27356
rect 24084 27344 24090 27396
rect 24578 27384 24584 27396
rect 24539 27356 24584 27384
rect 24578 27344 24584 27356
rect 24636 27344 24642 27396
rect 26326 27344 26332 27396
rect 26384 27384 26390 27396
rect 29089 27387 29147 27393
rect 29089 27384 29101 27387
rect 26384 27356 29101 27384
rect 26384 27344 26390 27356
rect 29089 27353 29101 27356
rect 29135 27353 29147 27387
rect 29089 27347 29147 27353
rect 29181 27387 29239 27393
rect 29181 27353 29193 27387
rect 29227 27384 29239 27387
rect 30466 27384 30472 27396
rect 29227 27356 30472 27384
rect 29227 27353 29239 27356
rect 29181 27347 29239 27353
rect 30466 27344 30472 27356
rect 30524 27344 30530 27396
rect 12066 27316 12072 27328
rect 7340 27288 7512 27316
rect 12027 27288 12072 27316
rect 7340 27276 7346 27288
rect 12066 27276 12072 27288
rect 12124 27316 12130 27328
rect 12342 27316 12348 27328
rect 12124 27288 12348 27316
rect 12124 27276 12130 27288
rect 12342 27276 12348 27288
rect 12400 27276 12406 27328
rect 19058 27325 19064 27328
rect 19015 27319 19064 27325
rect 19015 27285 19027 27319
rect 19061 27285 19064 27319
rect 19015 27279 19064 27285
rect 19058 27276 19064 27279
rect 19116 27276 19122 27328
rect 20162 27316 20168 27328
rect 20123 27288 20168 27316
rect 20162 27276 20168 27288
rect 20220 27276 20226 27328
rect 21913 27319 21971 27325
rect 21913 27285 21925 27319
rect 21959 27316 21971 27319
rect 22646 27316 22652 27328
rect 21959 27288 22652 27316
rect 21959 27285 21971 27288
rect 21913 27279 21971 27285
rect 22646 27276 22652 27288
rect 22704 27276 22710 27328
rect 22738 27276 22744 27328
rect 22796 27316 22802 27328
rect 22833 27319 22891 27325
rect 22833 27316 22845 27319
rect 22796 27288 22845 27316
rect 22796 27276 22802 27288
rect 22833 27285 22845 27288
rect 22879 27285 22891 27319
rect 30558 27316 30564 27328
rect 30519 27288 30564 27316
rect 22833 27279 22891 27285
rect 30558 27276 30564 27288
rect 30616 27276 30622 27328
rect 31202 27276 31208 27328
rect 31260 27316 31266 27328
rect 32401 27319 32459 27325
rect 32401 27316 32413 27319
rect 31260 27288 32413 27316
rect 31260 27276 31266 27288
rect 32401 27285 32413 27288
rect 32447 27285 32459 27319
rect 32582 27316 32588 27328
rect 32543 27288 32588 27316
rect 32401 27279 32459 27285
rect 32582 27276 32588 27288
rect 32640 27276 32646 27328
rect 1104 27226 34316 27248
rect 1104 27174 6517 27226
rect 6569 27174 6581 27226
rect 6633 27174 6645 27226
rect 6697 27174 6709 27226
rect 6761 27174 17588 27226
rect 17640 27174 17652 27226
rect 17704 27174 17716 27226
rect 17768 27174 17780 27226
rect 17832 27174 28658 27226
rect 28710 27174 28722 27226
rect 28774 27174 28786 27226
rect 28838 27174 28850 27226
rect 28902 27174 34316 27226
rect 1104 27152 34316 27174
rect 9858 27072 9864 27124
rect 9916 27112 9922 27124
rect 10413 27115 10471 27121
rect 10413 27112 10425 27115
rect 9916 27084 10425 27112
rect 9916 27072 9922 27084
rect 10413 27081 10425 27084
rect 10459 27081 10471 27115
rect 10413 27075 10471 27081
rect 11514 27072 11520 27124
rect 11572 27112 11578 27124
rect 12342 27112 12348 27124
rect 11572 27084 12348 27112
rect 11572 27072 11578 27084
rect 12342 27072 12348 27084
rect 12400 27072 12406 27124
rect 13446 27112 13452 27124
rect 13407 27084 13452 27112
rect 13446 27072 13452 27084
rect 13504 27072 13510 27124
rect 13538 27072 13544 27124
rect 13596 27112 13602 27124
rect 14645 27115 14703 27121
rect 14645 27112 14657 27115
rect 13596 27084 14657 27112
rect 13596 27072 13602 27084
rect 14645 27081 14657 27084
rect 14691 27081 14703 27115
rect 20162 27112 20168 27124
rect 14645 27075 14703 27081
rect 14844 27084 20168 27112
rect 11238 27004 11244 27056
rect 11296 27044 11302 27056
rect 13078 27044 13084 27056
rect 11296 27016 13084 27044
rect 11296 27004 11302 27016
rect 13078 27004 13084 27016
rect 13136 27044 13142 27056
rect 13357 27047 13415 27053
rect 13357 27044 13369 27047
rect 13136 27016 13369 27044
rect 13136 27004 13142 27016
rect 13357 27013 13369 27016
rect 13403 27044 13415 27047
rect 14093 27047 14151 27053
rect 14093 27044 14105 27047
rect 13403 27016 14105 27044
rect 13403 27013 13415 27016
rect 13357 27007 13415 27013
rect 14093 27013 14105 27016
rect 14139 27013 14151 27047
rect 14093 27007 14151 27013
rect 1486 26976 1492 26988
rect 1399 26948 1492 26976
rect 1486 26936 1492 26948
rect 1544 26976 1550 26988
rect 3973 26979 4031 26985
rect 1544 26948 1624 26976
rect 1544 26936 1550 26948
rect 1596 26908 1624 26948
rect 3973 26945 3985 26979
rect 4019 26976 4031 26979
rect 4019 26948 4660 26976
rect 4019 26945 4031 26948
rect 3973 26939 4031 26945
rect 1756 26911 1814 26917
rect 1596 26880 1716 26908
rect 1688 26840 1716 26880
rect 1756 26877 1768 26911
rect 1802 26908 1814 26911
rect 2682 26908 2688 26920
rect 1802 26880 2688 26908
rect 1802 26877 1814 26880
rect 1756 26871 1814 26877
rect 2682 26868 2688 26880
rect 2740 26868 2746 26920
rect 4522 26908 4528 26920
rect 2792 26880 4528 26908
rect 2792 26840 2820 26880
rect 4522 26868 4528 26880
rect 4580 26868 4586 26920
rect 4632 26908 4660 26948
rect 6086 26936 6092 26988
rect 6144 26976 6150 26988
rect 7926 26976 7932 26988
rect 6144 26948 7932 26976
rect 6144 26936 6150 26948
rect 7926 26936 7932 26948
rect 7984 26936 7990 26988
rect 8113 26979 8171 26985
rect 8113 26945 8125 26979
rect 8159 26976 8171 26979
rect 9030 26976 9036 26988
rect 8159 26948 9036 26976
rect 8159 26945 8171 26948
rect 8113 26939 8171 26945
rect 9030 26936 9036 26948
rect 9088 26936 9094 26988
rect 13446 26976 13452 26988
rect 12912 26948 13452 26976
rect 12912 26920 12940 26948
rect 13446 26936 13452 26948
rect 13504 26936 13510 26988
rect 13541 26979 13599 26985
rect 13541 26945 13553 26979
rect 13587 26976 13599 26979
rect 14182 26976 14188 26988
rect 13587 26948 14188 26976
rect 13587 26945 13599 26948
rect 13541 26939 13599 26945
rect 14182 26936 14188 26948
rect 14240 26936 14246 26988
rect 7837 26911 7895 26917
rect 4632 26880 5028 26908
rect 5000 26852 5028 26880
rect 7837 26877 7849 26911
rect 7883 26908 7895 26911
rect 8202 26908 8208 26920
rect 7883 26880 8208 26908
rect 7883 26877 7895 26880
rect 7837 26871 7895 26877
rect 8202 26868 8208 26880
rect 8260 26868 8266 26920
rect 8662 26908 8668 26920
rect 8623 26880 8668 26908
rect 8662 26868 8668 26880
rect 8720 26868 8726 26920
rect 8938 26908 8944 26920
rect 8899 26880 8944 26908
rect 8938 26868 8944 26880
rect 8996 26868 9002 26920
rect 9490 26908 9496 26920
rect 9451 26880 9496 26908
rect 9490 26868 9496 26880
rect 9548 26868 9554 26920
rect 10594 26908 10600 26920
rect 10555 26880 10600 26908
rect 10594 26868 10600 26880
rect 10652 26868 10658 26920
rect 10873 26911 10931 26917
rect 10873 26877 10885 26911
rect 10919 26908 10931 26911
rect 11146 26908 11152 26920
rect 10919 26880 11152 26908
rect 10919 26877 10931 26880
rect 10873 26871 10931 26877
rect 11146 26868 11152 26880
rect 11204 26868 11210 26920
rect 12434 26868 12440 26920
rect 12492 26908 12498 26920
rect 12894 26908 12900 26920
rect 12492 26880 12585 26908
rect 12855 26880 12900 26908
rect 12492 26868 12498 26880
rect 12894 26868 12900 26880
rect 12952 26868 12958 26920
rect 13262 26908 13268 26920
rect 13223 26880 13268 26908
rect 13262 26868 13268 26880
rect 13320 26868 13326 26920
rect 13814 26868 13820 26920
rect 13872 26908 13878 26920
rect 14844 26917 14872 27084
rect 20162 27072 20168 27084
rect 20220 27072 20226 27124
rect 22186 27072 22192 27124
rect 22244 27112 22250 27124
rect 22830 27112 22836 27124
rect 22244 27084 22836 27112
rect 22244 27072 22250 27084
rect 22830 27072 22836 27084
rect 22888 27112 22894 27124
rect 24762 27112 24768 27124
rect 22888 27084 23612 27112
rect 24723 27084 24768 27112
rect 22888 27072 22894 27084
rect 16393 27047 16451 27053
rect 16393 27013 16405 27047
rect 16439 27013 16451 27047
rect 16393 27007 16451 27013
rect 17589 27047 17647 27053
rect 17589 27013 17601 27047
rect 17635 27044 17647 27047
rect 22922 27044 22928 27056
rect 17635 27016 22928 27044
rect 17635 27013 17647 27016
rect 17589 27007 17647 27013
rect 16408 26976 16436 27007
rect 22922 27004 22928 27016
rect 22980 27004 22986 27056
rect 16666 26976 16672 26988
rect 16408 26948 16672 26976
rect 16666 26936 16672 26948
rect 16724 26976 16730 26988
rect 17954 26976 17960 26988
rect 16724 26948 17960 26976
rect 16724 26936 16730 26948
rect 17954 26936 17960 26948
rect 18012 26976 18018 26988
rect 18141 26979 18199 26985
rect 18141 26976 18153 26979
rect 18012 26948 18153 26976
rect 18012 26936 18018 26948
rect 18141 26945 18153 26948
rect 18187 26945 18199 26979
rect 19426 26976 19432 26988
rect 19387 26948 19432 26976
rect 18141 26939 18199 26945
rect 19426 26936 19432 26948
rect 19484 26936 19490 26988
rect 20714 26936 20720 26988
rect 20772 26976 20778 26988
rect 20901 26979 20959 26985
rect 20901 26976 20913 26979
rect 20772 26948 20913 26976
rect 20772 26936 20778 26948
rect 20901 26945 20913 26948
rect 20947 26945 20959 26979
rect 20901 26939 20959 26945
rect 21085 26979 21143 26985
rect 21085 26945 21097 26979
rect 21131 26976 21143 26979
rect 21174 26976 21180 26988
rect 21131 26948 21180 26976
rect 21131 26945 21143 26948
rect 21085 26939 21143 26945
rect 21174 26936 21180 26948
rect 21232 26936 21238 26988
rect 22738 26976 22744 26988
rect 22699 26948 22744 26976
rect 22738 26936 22744 26948
rect 22796 26936 22802 26988
rect 14001 26911 14059 26917
rect 14001 26908 14013 26911
rect 13872 26880 14013 26908
rect 13872 26868 13878 26880
rect 14001 26877 14013 26880
rect 14047 26877 14059 26911
rect 14001 26871 14059 26877
rect 14829 26911 14887 26917
rect 14829 26877 14841 26911
rect 14875 26877 14887 26911
rect 14829 26871 14887 26877
rect 14918 26868 14924 26920
rect 14976 26908 14982 26920
rect 15013 26911 15071 26917
rect 15013 26908 15025 26911
rect 14976 26880 15025 26908
rect 14976 26868 14982 26880
rect 15013 26877 15025 26880
rect 15059 26877 15071 26911
rect 15013 26871 15071 26877
rect 15280 26911 15338 26917
rect 15280 26877 15292 26911
rect 15326 26908 15338 26911
rect 16574 26908 16580 26920
rect 15326 26880 16580 26908
rect 15326 26877 15338 26880
rect 15280 26871 15338 26877
rect 16574 26868 16580 26880
rect 16632 26868 16638 26920
rect 17310 26908 17316 26920
rect 17271 26880 17316 26908
rect 17310 26868 17316 26880
rect 17368 26868 17374 26920
rect 17865 26911 17923 26917
rect 17865 26877 17877 26911
rect 17911 26877 17923 26911
rect 17865 26871 17923 26877
rect 3789 26843 3847 26849
rect 3789 26840 3801 26843
rect 1688 26812 2820 26840
rect 2884 26812 3801 26840
rect 2884 26784 2912 26812
rect 3789 26809 3801 26812
rect 3835 26809 3847 26843
rect 3789 26803 3847 26809
rect 4792 26843 4850 26849
rect 4792 26809 4804 26843
rect 4838 26840 4850 26843
rect 4890 26840 4896 26852
rect 4838 26812 4896 26840
rect 4838 26809 4850 26812
rect 4792 26803 4850 26809
rect 4890 26800 4896 26812
rect 4948 26800 4954 26852
rect 4982 26800 4988 26852
rect 5040 26800 5046 26852
rect 10318 26840 10324 26852
rect 5736 26812 10324 26840
rect 2866 26772 2872 26784
rect 2827 26744 2872 26772
rect 2866 26732 2872 26744
rect 2924 26732 2930 26784
rect 3326 26772 3332 26784
rect 3287 26744 3332 26772
rect 3326 26732 3332 26744
rect 3384 26732 3390 26784
rect 3697 26775 3755 26781
rect 3697 26741 3709 26775
rect 3743 26772 3755 26775
rect 5736 26772 5764 26812
rect 10318 26800 10324 26812
rect 10376 26800 10382 26852
rect 10781 26843 10839 26849
rect 10781 26809 10793 26843
rect 10827 26840 10839 26843
rect 12066 26840 12072 26852
rect 10827 26812 12072 26840
rect 10827 26809 10839 26812
rect 10781 26803 10839 26809
rect 12066 26800 12072 26812
rect 12124 26800 12130 26852
rect 12452 26840 12480 26868
rect 13280 26840 13308 26868
rect 12452 26812 13308 26840
rect 16592 26840 16620 26868
rect 17880 26840 17908 26871
rect 18598 26868 18604 26920
rect 18656 26908 18662 26920
rect 18969 26911 19027 26917
rect 18969 26908 18981 26911
rect 18656 26880 18981 26908
rect 18656 26868 18662 26880
rect 18969 26877 18981 26880
rect 19015 26877 19027 26911
rect 18969 26871 19027 26877
rect 19058 26868 19064 26920
rect 19116 26908 19122 26920
rect 20809 26911 20867 26917
rect 20809 26908 20821 26911
rect 19116 26880 20821 26908
rect 19116 26868 19122 26880
rect 20809 26877 20821 26880
rect 20855 26877 20867 26911
rect 20809 26871 20867 26877
rect 22186 26868 22192 26920
rect 22244 26908 22250 26920
rect 22557 26911 22615 26917
rect 22557 26908 22569 26911
rect 22244 26880 22569 26908
rect 22244 26868 22250 26880
rect 22557 26877 22569 26880
rect 22603 26877 22615 26911
rect 22557 26871 22615 26877
rect 22646 26868 22652 26920
rect 22704 26908 22710 26920
rect 22925 26911 22983 26917
rect 22704 26880 22749 26908
rect 22704 26868 22710 26880
rect 22925 26877 22937 26911
rect 22971 26877 22983 26911
rect 22925 26871 22983 26877
rect 22940 26840 22968 26871
rect 23014 26868 23020 26920
rect 23072 26908 23078 26920
rect 23584 26917 23612 27084
rect 24762 27072 24768 27084
rect 24820 27072 24826 27124
rect 31754 27112 31760 27124
rect 30760 27084 31760 27112
rect 24213 27047 24271 27053
rect 24213 27013 24225 27047
rect 24259 27044 24271 27047
rect 25038 27044 25044 27056
rect 24259 27016 25044 27044
rect 24259 27013 24271 27016
rect 24213 27007 24271 27013
rect 25038 27004 25044 27016
rect 25096 27004 25102 27056
rect 27614 27004 27620 27056
rect 27672 27044 27678 27056
rect 30760 27044 30788 27084
rect 31754 27072 31760 27084
rect 31812 27072 31818 27124
rect 27672 27016 30788 27044
rect 27672 27004 27678 27016
rect 25314 26936 25320 26988
rect 25372 26976 25378 26988
rect 27893 26979 27951 26985
rect 27893 26976 27905 26979
rect 25372 26948 27905 26976
rect 25372 26936 25378 26948
rect 27893 26945 27905 26948
rect 27939 26945 27951 26979
rect 29822 26976 29828 26988
rect 29783 26948 29828 26976
rect 27893 26939 27951 26945
rect 29822 26936 29828 26948
rect 29880 26936 29886 26988
rect 30760 26985 30788 27016
rect 30745 26979 30803 26985
rect 30745 26945 30757 26979
rect 30791 26945 30803 26979
rect 33226 26976 33232 26988
rect 30745 26939 30803 26945
rect 33060 26948 33232 26976
rect 23385 26911 23443 26917
rect 23385 26908 23397 26911
rect 23072 26880 23397 26908
rect 23072 26868 23078 26880
rect 23385 26877 23397 26880
rect 23431 26877 23443 26911
rect 23385 26871 23443 26877
rect 23569 26911 23627 26917
rect 23569 26877 23581 26911
rect 23615 26877 23627 26911
rect 24026 26908 24032 26920
rect 23987 26880 24032 26908
rect 23569 26871 23627 26877
rect 24026 26868 24032 26880
rect 24084 26868 24090 26920
rect 24305 26911 24363 26917
rect 24305 26877 24317 26911
rect 24351 26877 24363 26911
rect 24305 26871 24363 26877
rect 24581 26911 24639 26917
rect 24581 26877 24593 26911
rect 24627 26908 24639 26911
rect 26234 26908 26240 26920
rect 24627 26880 26240 26908
rect 24627 26877 24639 26880
rect 24581 26871 24639 26877
rect 23477 26843 23535 26849
rect 23477 26840 23489 26843
rect 16592 26812 17908 26840
rect 22066 26812 22876 26840
rect 22940 26812 23489 26840
rect 5902 26772 5908 26784
rect 3743 26744 5764 26772
rect 5863 26744 5908 26772
rect 3743 26741 3755 26744
rect 3697 26735 3755 26741
rect 5902 26732 5908 26744
rect 5960 26732 5966 26784
rect 7466 26772 7472 26784
rect 7427 26744 7472 26772
rect 7466 26732 7472 26744
rect 7524 26732 7530 26784
rect 8754 26772 8760 26784
rect 8715 26744 8760 26772
rect 8754 26732 8760 26744
rect 8812 26732 8818 26784
rect 13081 26775 13139 26781
rect 13081 26741 13093 26775
rect 13127 26772 13139 26775
rect 13630 26772 13636 26784
rect 13127 26744 13636 26772
rect 13127 26741 13139 26744
rect 13081 26735 13139 26741
rect 13630 26732 13636 26744
rect 13688 26732 13694 26784
rect 20438 26772 20444 26784
rect 20399 26744 20444 26772
rect 20438 26732 20444 26744
rect 20496 26732 20502 26784
rect 21082 26732 21088 26784
rect 21140 26772 21146 26784
rect 22066 26772 22094 26812
rect 22848 26781 22876 26812
rect 23477 26809 23489 26812
rect 23523 26809 23535 26843
rect 24320 26840 24348 26871
rect 26234 26868 26240 26880
rect 26292 26868 26298 26920
rect 27798 26868 27804 26920
rect 27856 26908 27862 26920
rect 27985 26911 28043 26917
rect 27985 26908 27997 26911
rect 27856 26880 27997 26908
rect 27856 26868 27862 26880
rect 27985 26877 27997 26880
rect 28031 26877 28043 26911
rect 30098 26908 30104 26920
rect 30059 26880 30104 26908
rect 27985 26871 28043 26877
rect 30098 26868 30104 26880
rect 30156 26868 30162 26920
rect 31012 26911 31070 26917
rect 31012 26877 31024 26911
rect 31058 26908 31070 26911
rect 33060 26908 33088 26948
rect 33226 26936 33232 26948
rect 33284 26976 33290 26988
rect 33284 26948 33364 26976
rect 33284 26936 33290 26948
rect 33336 26917 33364 26948
rect 31058 26880 33088 26908
rect 33137 26911 33195 26917
rect 31058 26877 31070 26880
rect 31012 26871 31070 26877
rect 33137 26877 33149 26911
rect 33183 26877 33195 26911
rect 33137 26871 33195 26877
rect 33321 26911 33379 26917
rect 33321 26877 33333 26911
rect 33367 26877 33379 26911
rect 33321 26871 33379 26877
rect 24854 26840 24860 26852
rect 24320 26812 24860 26840
rect 23477 26803 23535 26809
rect 24854 26800 24860 26812
rect 24912 26800 24918 26852
rect 31570 26800 31576 26852
rect 31628 26840 31634 26852
rect 33045 26843 33103 26849
rect 33045 26840 33057 26843
rect 31628 26812 33057 26840
rect 31628 26800 31634 26812
rect 33045 26809 33057 26812
rect 33091 26809 33103 26843
rect 33045 26803 33103 26809
rect 21140 26744 22094 26772
rect 22833 26775 22891 26781
rect 21140 26732 21146 26744
rect 22833 26741 22845 26775
rect 22879 26741 22891 26775
rect 22833 26735 22891 26741
rect 24397 26775 24455 26781
rect 24397 26741 24409 26775
rect 24443 26772 24455 26775
rect 24946 26772 24952 26784
rect 24443 26744 24952 26772
rect 24443 26741 24455 26744
rect 24397 26735 24455 26741
rect 24946 26732 24952 26744
rect 25004 26732 25010 26784
rect 28166 26732 28172 26784
rect 28224 26772 28230 26784
rect 28353 26775 28411 26781
rect 28353 26772 28365 26775
rect 28224 26744 28365 26772
rect 28224 26732 28230 26744
rect 28353 26741 28365 26744
rect 28399 26741 28411 26775
rect 28353 26735 28411 26741
rect 32125 26775 32183 26781
rect 32125 26741 32137 26775
rect 32171 26772 32183 26775
rect 32950 26772 32956 26784
rect 32171 26744 32956 26772
rect 32171 26741 32183 26744
rect 32125 26735 32183 26741
rect 32950 26732 32956 26744
rect 33008 26772 33014 26784
rect 33152 26772 33180 26871
rect 33008 26744 33180 26772
rect 33008 26732 33014 26744
rect 1104 26682 34316 26704
rect 1104 26630 12052 26682
rect 12104 26630 12116 26682
rect 12168 26630 12180 26682
rect 12232 26630 12244 26682
rect 12296 26630 23123 26682
rect 23175 26630 23187 26682
rect 23239 26630 23251 26682
rect 23303 26630 23315 26682
rect 23367 26630 34316 26682
rect 1104 26608 34316 26630
rect 2961 26571 3019 26577
rect 2961 26537 2973 26571
rect 3007 26568 3019 26571
rect 3142 26568 3148 26580
rect 3007 26540 3148 26568
rect 3007 26537 3019 26540
rect 2961 26531 3019 26537
rect 3142 26528 3148 26540
rect 3200 26528 3206 26580
rect 4890 26568 4896 26580
rect 4851 26540 4896 26568
rect 4890 26528 4896 26540
rect 4948 26528 4954 26580
rect 7466 26568 7472 26580
rect 7427 26540 7472 26568
rect 7466 26528 7472 26540
rect 7524 26528 7530 26580
rect 8386 26568 8392 26580
rect 8347 26540 8392 26568
rect 8386 26528 8392 26540
rect 8444 26528 8450 26580
rect 10045 26571 10103 26577
rect 10045 26537 10057 26571
rect 10091 26568 10103 26571
rect 10226 26568 10232 26580
rect 10091 26540 10232 26568
rect 10091 26537 10103 26540
rect 10045 26531 10103 26537
rect 10226 26528 10232 26540
rect 10284 26528 10290 26580
rect 16574 26528 16580 26580
rect 16632 26568 16638 26580
rect 16761 26571 16819 26577
rect 16761 26568 16773 26571
rect 16632 26540 16773 26568
rect 16632 26528 16638 26540
rect 16761 26537 16773 26540
rect 16807 26537 16819 26571
rect 16761 26531 16819 26537
rect 18966 26528 18972 26580
rect 19024 26568 19030 26580
rect 19061 26571 19119 26577
rect 19061 26568 19073 26571
rect 19024 26540 19073 26568
rect 19024 26528 19030 26540
rect 19061 26537 19073 26540
rect 19107 26537 19119 26571
rect 19061 26531 19119 26537
rect 19426 26528 19432 26580
rect 19484 26568 19490 26580
rect 20162 26568 20168 26580
rect 19484 26540 20168 26568
rect 19484 26528 19490 26540
rect 20162 26528 20168 26540
rect 20220 26568 20226 26580
rect 20220 26540 21496 26568
rect 20220 26528 20226 26540
rect 1578 26460 1584 26512
rect 1636 26500 1642 26512
rect 7377 26503 7435 26509
rect 7377 26500 7389 26503
rect 1636 26472 7389 26500
rect 1636 26460 1642 26472
rect 7377 26469 7389 26472
rect 7423 26469 7435 26503
rect 7377 26463 7435 26469
rect 10134 26460 10140 26512
rect 10192 26500 10198 26512
rect 11333 26503 11391 26509
rect 11333 26500 11345 26503
rect 10192 26472 11345 26500
rect 10192 26460 10198 26472
rect 11333 26469 11345 26472
rect 11379 26469 11391 26503
rect 11333 26463 11391 26469
rect 12158 26460 12164 26512
rect 12216 26500 12222 26512
rect 12253 26503 12311 26509
rect 12253 26500 12265 26503
rect 12216 26472 12265 26500
rect 12216 26460 12222 26472
rect 12253 26469 12265 26472
rect 12299 26469 12311 26503
rect 12253 26463 12311 26469
rect 12434 26460 12440 26512
rect 12492 26509 12498 26512
rect 12492 26503 12516 26509
rect 12504 26469 12516 26503
rect 12492 26463 12516 26469
rect 13449 26503 13507 26509
rect 13449 26469 13461 26503
rect 13495 26500 13507 26503
rect 13541 26503 13599 26509
rect 13541 26500 13553 26503
rect 13495 26472 13553 26500
rect 13495 26469 13507 26472
rect 13449 26463 13507 26469
rect 13541 26469 13553 26472
rect 13587 26500 13599 26503
rect 13814 26500 13820 26512
rect 13587 26472 13820 26500
rect 13587 26469 13599 26472
rect 13541 26463 13599 26469
rect 12492 26460 12498 26463
rect 13814 26460 13820 26472
rect 13872 26460 13878 26512
rect 14734 26500 14740 26512
rect 14695 26472 14740 26500
rect 14734 26460 14740 26472
rect 14792 26460 14798 26512
rect 16666 26500 16672 26512
rect 16627 26472 16672 26500
rect 16666 26460 16672 26472
rect 16724 26460 16730 26512
rect 21468 26486 21496 26540
rect 22922 26528 22928 26580
rect 22980 26568 22986 26580
rect 25314 26568 25320 26580
rect 22980 26540 25320 26568
rect 22980 26528 22986 26540
rect 25314 26528 25320 26540
rect 25372 26528 25378 26580
rect 27798 26568 27804 26580
rect 27759 26540 27804 26568
rect 27798 26528 27804 26540
rect 27856 26528 27862 26580
rect 33137 26571 33195 26577
rect 33137 26537 33149 26571
rect 33183 26568 33195 26571
rect 33226 26568 33232 26580
rect 33183 26540 33232 26568
rect 33183 26537 33195 26540
rect 33137 26531 33195 26537
rect 33226 26528 33232 26540
rect 33284 26528 33290 26580
rect 22511 26503 22569 26509
rect 22511 26469 22523 26503
rect 22557 26500 22569 26503
rect 23014 26500 23020 26512
rect 22557 26472 23020 26500
rect 22557 26469 22569 26472
rect 22511 26463 22569 26469
rect 23014 26460 23020 26472
rect 23072 26500 23078 26512
rect 26326 26500 26332 26512
rect 23072 26472 23336 26500
rect 26287 26472 26332 26500
rect 23072 26460 23078 26472
rect 2866 26392 2872 26444
rect 2924 26432 2930 26444
rect 3145 26435 3203 26441
rect 3145 26432 3157 26435
rect 2924 26404 3157 26432
rect 2924 26392 2930 26404
rect 3145 26401 3157 26404
rect 3191 26401 3203 26435
rect 3145 26395 3203 26401
rect 4430 26392 4436 26444
rect 4488 26432 4494 26444
rect 5074 26432 5080 26444
rect 4488 26404 5080 26432
rect 4488 26392 4494 26404
rect 5074 26392 5080 26404
rect 5132 26392 5138 26444
rect 5169 26435 5227 26441
rect 5169 26401 5181 26435
rect 5215 26432 5227 26435
rect 5902 26432 5908 26444
rect 5215 26404 5908 26432
rect 5215 26401 5227 26404
rect 5169 26395 5227 26401
rect 5902 26392 5908 26404
rect 5960 26392 5966 26444
rect 7926 26392 7932 26444
rect 7984 26432 7990 26444
rect 8297 26435 8355 26441
rect 8297 26432 8309 26435
rect 7984 26404 8309 26432
rect 7984 26392 7990 26404
rect 8297 26401 8309 26404
rect 8343 26401 8355 26435
rect 10410 26432 10416 26444
rect 10371 26404 10416 26432
rect 8297 26395 8355 26401
rect 10410 26392 10416 26404
rect 10468 26392 10474 26444
rect 10594 26392 10600 26444
rect 10652 26432 10658 26444
rect 10652 26404 10732 26432
rect 10652 26392 10658 26404
rect 3329 26367 3387 26373
rect 3329 26333 3341 26367
rect 3375 26364 3387 26367
rect 4338 26364 4344 26376
rect 3375 26336 4344 26364
rect 3375 26333 3387 26336
rect 3329 26327 3387 26333
rect 4338 26324 4344 26336
rect 4396 26324 4402 26376
rect 5534 26364 5540 26376
rect 5495 26336 5540 26364
rect 5534 26324 5540 26336
rect 5592 26324 5598 26376
rect 7190 26364 7196 26376
rect 7151 26336 7196 26364
rect 7190 26324 7196 26336
rect 7248 26324 7254 26376
rect 10704 26373 10732 26404
rect 10870 26392 10876 26444
rect 10928 26432 10934 26444
rect 11609 26435 11667 26441
rect 11609 26432 11621 26435
rect 10928 26404 11621 26432
rect 10928 26392 10934 26404
rect 11609 26401 11621 26404
rect 11655 26432 11667 26435
rect 11974 26432 11980 26444
rect 11655 26404 11980 26432
rect 11655 26401 11667 26404
rect 11609 26395 11667 26401
rect 11974 26392 11980 26404
rect 12032 26392 12038 26444
rect 13725 26435 13783 26441
rect 13725 26401 13737 26435
rect 13771 26432 13783 26435
rect 14550 26432 14556 26444
rect 13771 26404 14556 26432
rect 13771 26401 13783 26404
rect 13725 26395 13783 26401
rect 14550 26392 14556 26404
rect 14608 26432 14614 26444
rect 14921 26435 14979 26441
rect 14921 26432 14933 26435
rect 14608 26404 14933 26432
rect 14608 26392 14614 26404
rect 14921 26401 14933 26404
rect 14967 26401 14979 26435
rect 15562 26432 15568 26444
rect 15523 26404 15568 26432
rect 14921 26395 14979 26401
rect 15562 26392 15568 26404
rect 15620 26392 15626 26444
rect 16945 26435 17003 26441
rect 16945 26401 16957 26435
rect 16991 26432 17003 26435
rect 17310 26432 17316 26444
rect 16991 26404 17316 26432
rect 16991 26401 17003 26404
rect 16945 26395 17003 26401
rect 17310 26392 17316 26404
rect 17368 26392 17374 26444
rect 18690 26432 18696 26444
rect 18651 26404 18696 26432
rect 18690 26392 18696 26404
rect 18748 26392 18754 26444
rect 18877 26435 18935 26441
rect 18877 26401 18889 26435
rect 18923 26432 18935 26435
rect 19058 26432 19064 26444
rect 18923 26404 19064 26432
rect 18923 26401 18935 26404
rect 18877 26395 18935 26401
rect 19058 26392 19064 26404
rect 19116 26392 19122 26444
rect 21082 26432 21088 26444
rect 21043 26404 21088 26432
rect 21082 26392 21088 26404
rect 21140 26392 21146 26444
rect 22278 26392 22284 26444
rect 22336 26432 22342 26444
rect 23308 26441 23336 26472
rect 26326 26460 26332 26472
rect 26384 26460 26390 26512
rect 30098 26500 30104 26512
rect 27554 26472 30104 26500
rect 30098 26460 30104 26472
rect 30156 26460 30162 26512
rect 33502 26500 33508 26512
rect 30944 26472 33508 26500
rect 23109 26435 23167 26441
rect 23109 26432 23121 26435
rect 22336 26404 23121 26432
rect 22336 26392 22342 26404
rect 23109 26401 23121 26404
rect 23155 26401 23167 26435
rect 23109 26395 23167 26401
rect 23293 26435 23351 26441
rect 23293 26401 23305 26435
rect 23339 26401 23351 26435
rect 23293 26395 23351 26401
rect 24121 26435 24179 26441
rect 24121 26401 24133 26435
rect 24167 26401 24179 26435
rect 24121 26395 24179 26401
rect 24305 26435 24363 26441
rect 24305 26401 24317 26435
rect 24351 26401 24363 26435
rect 25314 26432 25320 26444
rect 25275 26404 25320 26432
rect 24305 26395 24363 26401
rect 10505 26367 10563 26373
rect 10505 26333 10517 26367
rect 10551 26364 10563 26367
rect 10689 26367 10747 26373
rect 10551 26336 10640 26364
rect 10551 26333 10563 26336
rect 10505 26327 10563 26333
rect 7834 26228 7840 26240
rect 7795 26200 7840 26228
rect 7834 26188 7840 26200
rect 7892 26188 7898 26240
rect 9030 26188 9036 26240
rect 9088 26228 9094 26240
rect 10612 26228 10640 26336
rect 10689 26333 10701 26367
rect 10735 26333 10747 26367
rect 11238 26364 11244 26376
rect 11199 26336 11244 26364
rect 10689 26327 10747 26333
rect 10704 26296 10732 26327
rect 11238 26324 11244 26336
rect 11296 26324 11302 26376
rect 11422 26324 11428 26376
rect 11480 26364 11486 26376
rect 11793 26367 11851 26373
rect 11793 26364 11805 26367
rect 11480 26336 11805 26364
rect 11480 26324 11486 26336
rect 11793 26333 11805 26336
rect 11839 26333 11851 26367
rect 15580 26364 15608 26392
rect 11793 26327 11851 26333
rect 11900 26336 15608 26364
rect 20717 26367 20775 26373
rect 11900 26296 11928 26336
rect 20717 26333 20729 26367
rect 20763 26364 20775 26367
rect 20898 26364 20904 26376
rect 20763 26336 20904 26364
rect 20763 26333 20775 26336
rect 20717 26327 20775 26333
rect 20898 26324 20904 26336
rect 20956 26324 20962 26376
rect 22370 26324 22376 26376
rect 22428 26364 22434 26376
rect 23017 26367 23075 26373
rect 23017 26364 23029 26367
rect 22428 26336 23029 26364
rect 22428 26324 22434 26336
rect 23017 26333 23029 26336
rect 23063 26333 23075 26367
rect 23124 26364 23152 26395
rect 23937 26367 23995 26373
rect 23937 26364 23949 26367
rect 23124 26336 23949 26364
rect 23017 26327 23075 26333
rect 23937 26333 23949 26336
rect 23983 26333 23995 26367
rect 23937 26327 23995 26333
rect 12802 26296 12808 26308
rect 10704 26268 11928 26296
rect 12452 26268 12808 26296
rect 11882 26228 11888 26240
rect 9088 26200 11888 26228
rect 9088 26188 9094 26200
rect 11882 26188 11888 26200
rect 11940 26188 11946 26240
rect 12452 26237 12480 26268
rect 12802 26256 12808 26268
rect 12860 26296 12866 26308
rect 13449 26299 13507 26305
rect 13449 26296 13461 26299
rect 12860 26268 13461 26296
rect 12860 26256 12866 26268
rect 13449 26265 13461 26268
rect 13495 26265 13507 26299
rect 13449 26259 13507 26265
rect 17129 26299 17187 26305
rect 17129 26265 17141 26299
rect 17175 26296 17187 26299
rect 18782 26296 18788 26308
rect 17175 26268 18788 26296
rect 17175 26265 17187 26268
rect 17129 26259 17187 26265
rect 18782 26256 18788 26268
rect 18840 26256 18846 26308
rect 24136 26296 24164 26395
rect 24320 26364 24348 26395
rect 25314 26392 25320 26404
rect 25372 26392 25378 26444
rect 25406 26392 25412 26444
rect 25464 26432 25470 26444
rect 30944 26441 30972 26472
rect 33502 26460 33508 26472
rect 33560 26460 33566 26512
rect 25501 26435 25559 26441
rect 25501 26432 25513 26435
rect 25464 26404 25513 26432
rect 25464 26392 25470 26404
rect 25501 26401 25513 26404
rect 25547 26401 25559 26435
rect 25501 26395 25559 26401
rect 29365 26435 29423 26441
rect 29365 26401 29377 26435
rect 29411 26401 29423 26435
rect 29365 26395 29423 26401
rect 29549 26435 29607 26441
rect 29549 26401 29561 26435
rect 29595 26432 29607 26435
rect 30929 26435 30987 26441
rect 30929 26432 30941 26435
rect 29595 26404 30941 26432
rect 29595 26401 29607 26404
rect 29549 26395 29607 26401
rect 30929 26401 30941 26404
rect 30975 26401 30987 26435
rect 31294 26432 31300 26444
rect 31255 26404 31300 26432
rect 30929 26395 30987 26401
rect 24854 26364 24860 26376
rect 24320 26336 24860 26364
rect 24854 26324 24860 26336
rect 24912 26364 24918 26376
rect 26053 26367 26111 26373
rect 24912 26336 25544 26364
rect 24912 26324 24918 26336
rect 25516 26308 25544 26336
rect 26053 26333 26065 26367
rect 26099 26364 26111 26367
rect 27614 26364 27620 26376
rect 26099 26336 27620 26364
rect 26099 26333 26111 26336
rect 26053 26327 26111 26333
rect 27614 26324 27620 26336
rect 27672 26324 27678 26376
rect 29380 26364 29408 26395
rect 31294 26392 31300 26404
rect 31352 26392 31358 26444
rect 32024 26435 32082 26441
rect 32024 26432 32036 26435
rect 31404 26404 32036 26432
rect 30558 26364 30564 26376
rect 29380 26336 30564 26364
rect 30558 26324 30564 26336
rect 30616 26364 30622 26376
rect 30745 26367 30803 26373
rect 30745 26364 30757 26367
rect 30616 26336 30757 26364
rect 30616 26324 30622 26336
rect 30745 26333 30757 26336
rect 30791 26364 30803 26367
rect 31404 26364 31432 26404
rect 32024 26401 32036 26404
rect 32070 26432 32082 26435
rect 32582 26432 32588 26444
rect 32070 26404 32588 26432
rect 32070 26401 32082 26404
rect 32024 26395 32082 26401
rect 32582 26392 32588 26404
rect 32640 26432 32646 26444
rect 33042 26432 33048 26444
rect 32640 26404 33048 26432
rect 32640 26392 32646 26404
rect 33042 26392 33048 26404
rect 33100 26392 33106 26444
rect 31754 26364 31760 26376
rect 30791 26336 31432 26364
rect 31715 26336 31760 26364
rect 30791 26333 30803 26336
rect 30745 26327 30803 26333
rect 31754 26324 31760 26336
rect 31812 26324 31818 26376
rect 24946 26296 24952 26308
rect 24136 26268 24952 26296
rect 24946 26256 24952 26268
rect 25004 26256 25010 26308
rect 25498 26296 25504 26308
rect 25459 26268 25504 26296
rect 25498 26256 25504 26268
rect 25556 26256 25562 26308
rect 31205 26299 31263 26305
rect 31205 26265 31217 26299
rect 31251 26296 31263 26299
rect 31251 26268 31800 26296
rect 31251 26265 31263 26268
rect 31205 26259 31263 26265
rect 31772 26240 31800 26268
rect 12437 26231 12495 26237
rect 12437 26197 12449 26231
rect 12483 26197 12495 26231
rect 12437 26191 12495 26197
rect 12618 26188 12624 26240
rect 12676 26228 12682 26240
rect 12676 26200 12721 26228
rect 12676 26188 12682 26200
rect 29362 26188 29368 26240
rect 29420 26228 29426 26240
rect 29457 26231 29515 26237
rect 29457 26228 29469 26231
rect 29420 26200 29469 26228
rect 29420 26188 29426 26200
rect 29457 26197 29469 26200
rect 29503 26197 29515 26231
rect 29457 26191 29515 26197
rect 31754 26188 31760 26240
rect 31812 26188 31818 26240
rect 1104 26138 34316 26160
rect 1104 26086 6517 26138
rect 6569 26086 6581 26138
rect 6633 26086 6645 26138
rect 6697 26086 6709 26138
rect 6761 26086 17588 26138
rect 17640 26086 17652 26138
rect 17704 26086 17716 26138
rect 17768 26086 17780 26138
rect 17832 26086 28658 26138
rect 28710 26086 28722 26138
rect 28774 26086 28786 26138
rect 28838 26086 28850 26138
rect 28902 26086 34316 26138
rect 1104 26064 34316 26086
rect 4893 26027 4951 26033
rect 4893 25993 4905 26027
rect 4939 26024 4951 26027
rect 5534 26024 5540 26036
rect 4939 25996 5540 26024
rect 4939 25993 4951 25996
rect 4893 25987 4951 25993
rect 5534 25984 5540 25996
rect 5592 25984 5598 26036
rect 7929 26027 7987 26033
rect 7929 25993 7941 26027
rect 7975 26024 7987 26027
rect 8662 26024 8668 26036
rect 7975 25996 8668 26024
rect 7975 25993 7987 25996
rect 7929 25987 7987 25993
rect 8662 25984 8668 25996
rect 8720 25984 8726 26036
rect 10410 25984 10416 26036
rect 10468 26024 10474 26036
rect 10505 26027 10563 26033
rect 10505 26024 10517 26027
rect 10468 25996 10517 26024
rect 10468 25984 10474 25996
rect 10505 25993 10517 25996
rect 10551 25993 10563 26027
rect 10505 25987 10563 25993
rect 12713 26027 12771 26033
rect 12713 25993 12725 26027
rect 12759 26024 12771 26027
rect 13814 26024 13820 26036
rect 12759 25996 13820 26024
rect 12759 25993 12771 25996
rect 12713 25987 12771 25993
rect 13814 25984 13820 25996
rect 13872 25984 13878 26036
rect 14550 26024 14556 26036
rect 14511 25996 14556 26024
rect 14550 25984 14556 25996
rect 14608 25984 14614 26036
rect 15010 25984 15016 26036
rect 15068 26024 15074 26036
rect 15068 25996 20392 26024
rect 15068 25984 15074 25996
rect 7190 25916 7196 25968
rect 7248 25956 7254 25968
rect 9766 25956 9772 25968
rect 7248 25928 9772 25956
rect 7248 25916 7254 25928
rect 9766 25916 9772 25928
rect 9824 25916 9830 25968
rect 10965 25959 11023 25965
rect 10965 25925 10977 25959
rect 11011 25925 11023 25959
rect 11146 25956 11152 25968
rect 10965 25919 11023 25925
rect 11072 25928 11152 25956
rect 3234 25848 3240 25900
rect 3292 25888 3298 25900
rect 3421 25891 3479 25897
rect 3421 25888 3433 25891
rect 3292 25860 3433 25888
rect 3292 25848 3298 25860
rect 3421 25857 3433 25860
rect 3467 25888 3479 25891
rect 7282 25888 7288 25900
rect 3467 25860 5488 25888
rect 7243 25860 7288 25888
rect 3467 25857 3479 25860
rect 3421 25851 3479 25857
rect 5074 25820 5080 25832
rect 5035 25792 5080 25820
rect 5074 25780 5080 25792
rect 5132 25780 5138 25832
rect 5258 25780 5264 25832
rect 5316 25820 5322 25832
rect 5353 25823 5411 25829
rect 5353 25820 5365 25823
rect 5316 25792 5365 25820
rect 5316 25780 5322 25792
rect 5353 25789 5365 25792
rect 5399 25789 5411 25823
rect 5353 25783 5411 25789
rect 2774 25712 2780 25764
rect 2832 25752 2838 25764
rect 3145 25755 3203 25761
rect 3145 25752 3157 25755
rect 2832 25724 3157 25752
rect 2832 25712 2838 25724
rect 3145 25721 3157 25724
rect 3191 25752 3203 25755
rect 5276 25752 5304 25780
rect 3191 25724 5304 25752
rect 3191 25721 3203 25724
rect 3145 25715 3203 25721
rect 4982 25644 4988 25696
rect 5040 25684 5046 25696
rect 5261 25687 5319 25693
rect 5261 25684 5273 25687
rect 5040 25656 5273 25684
rect 5040 25644 5046 25656
rect 5261 25653 5273 25656
rect 5307 25653 5319 25687
rect 5460 25684 5488 25860
rect 7282 25848 7288 25860
rect 7340 25848 7346 25900
rect 7466 25888 7472 25900
rect 7427 25860 7472 25888
rect 7466 25848 7472 25860
rect 7524 25848 7530 25900
rect 8941 25891 8999 25897
rect 8941 25857 8953 25891
rect 8987 25888 8999 25891
rect 9030 25888 9036 25900
rect 8987 25860 9036 25888
rect 8987 25857 8999 25860
rect 8941 25851 8999 25857
rect 9030 25848 9036 25860
rect 9088 25848 9094 25900
rect 10980 25888 11008 25919
rect 9140 25860 11008 25888
rect 7561 25823 7619 25829
rect 7561 25789 7573 25823
rect 7607 25820 7619 25823
rect 7834 25820 7840 25832
rect 7607 25792 7840 25820
rect 7607 25789 7619 25792
rect 7561 25783 7619 25789
rect 7834 25780 7840 25792
rect 7892 25780 7898 25832
rect 8754 25820 8760 25832
rect 7944 25792 8760 25820
rect 7374 25712 7380 25764
rect 7432 25752 7438 25764
rect 7944 25752 7972 25792
rect 8754 25780 8760 25792
rect 8812 25820 8818 25832
rect 9140 25820 9168 25860
rect 10318 25820 10324 25832
rect 8812 25792 9168 25820
rect 10279 25792 10324 25820
rect 8812 25780 8818 25792
rect 10318 25780 10324 25792
rect 10376 25780 10382 25832
rect 10505 25823 10563 25829
rect 10505 25789 10517 25823
rect 10551 25820 10563 25823
rect 11072 25820 11100 25928
rect 11146 25916 11152 25928
rect 11204 25916 11210 25968
rect 11422 25916 11428 25968
rect 11480 25956 11486 25968
rect 12161 25959 12219 25965
rect 12161 25956 12173 25959
rect 11480 25928 12173 25956
rect 11480 25916 11486 25928
rect 12161 25925 12173 25928
rect 12207 25956 12219 25959
rect 12434 25956 12440 25968
rect 12207 25928 12440 25956
rect 12207 25925 12219 25928
rect 12161 25919 12219 25925
rect 12434 25916 12440 25928
rect 12492 25916 12498 25968
rect 20364 25956 20392 25996
rect 20714 25984 20720 26036
rect 20772 26024 20778 26036
rect 21039 26027 21097 26033
rect 21039 26024 21051 26027
rect 20772 25996 21051 26024
rect 20772 25984 20778 25996
rect 21039 25993 21051 25996
rect 21085 25993 21097 26027
rect 21039 25987 21097 25993
rect 22462 25984 22468 26036
rect 22520 26024 22526 26036
rect 22833 26027 22891 26033
rect 22833 26024 22845 26027
rect 22520 25996 22845 26024
rect 22520 25984 22526 25996
rect 22833 25993 22845 25996
rect 22879 25993 22891 26027
rect 22833 25987 22891 25993
rect 26510 25984 26516 26036
rect 26568 26024 26574 26036
rect 27522 26024 27528 26036
rect 26568 25996 27528 26024
rect 26568 25984 26574 25996
rect 27522 25984 27528 25996
rect 27580 26024 27586 26036
rect 30374 26024 30380 26036
rect 27580 25996 30380 26024
rect 27580 25984 27586 25996
rect 30374 25984 30380 25996
rect 30432 25984 30438 26036
rect 30926 25956 30932 25968
rect 20364 25928 26924 25956
rect 30887 25928 30932 25956
rect 13630 25888 13636 25900
rect 11164 25860 13636 25888
rect 11164 25829 11192 25860
rect 13630 25848 13636 25860
rect 13688 25848 13694 25900
rect 19613 25891 19671 25897
rect 19613 25857 19625 25891
rect 19659 25888 19671 25891
rect 20438 25888 20444 25900
rect 19659 25860 20444 25888
rect 19659 25857 19671 25860
rect 19613 25851 19671 25857
rect 20438 25848 20444 25860
rect 20496 25848 20502 25900
rect 26326 25888 26332 25900
rect 25240 25860 26332 25888
rect 10551 25792 11100 25820
rect 11149 25823 11207 25829
rect 10551 25789 10563 25792
rect 10505 25783 10563 25789
rect 11149 25789 11161 25823
rect 11195 25789 11207 25823
rect 11149 25783 11207 25789
rect 11698 25780 11704 25832
rect 11756 25820 11762 25832
rect 12069 25823 12127 25829
rect 12069 25820 12081 25823
rect 11756 25792 12081 25820
rect 11756 25780 11762 25792
rect 12069 25789 12081 25792
rect 12115 25789 12127 25823
rect 12069 25783 12127 25789
rect 12253 25823 12311 25829
rect 12253 25789 12265 25823
rect 12299 25820 12311 25823
rect 12342 25820 12348 25832
rect 12299 25792 12348 25820
rect 12299 25789 12311 25792
rect 12253 25783 12311 25789
rect 7432 25724 7972 25752
rect 9125 25755 9183 25761
rect 7432 25712 7438 25724
rect 9125 25721 9137 25755
rect 9171 25752 9183 25755
rect 10778 25752 10784 25764
rect 9171 25724 10784 25752
rect 9171 25721 9183 25724
rect 9125 25715 9183 25721
rect 10778 25712 10784 25724
rect 10836 25712 10842 25764
rect 11790 25712 11796 25764
rect 11848 25752 11854 25764
rect 12268 25752 12296 25783
rect 12342 25780 12348 25792
rect 12400 25780 12406 25832
rect 12713 25823 12771 25829
rect 12713 25789 12725 25823
rect 12759 25820 12771 25823
rect 12805 25823 12863 25829
rect 12805 25820 12817 25823
rect 12759 25792 12817 25820
rect 12759 25789 12771 25792
rect 12713 25783 12771 25789
rect 12805 25789 12817 25792
rect 12851 25789 12863 25823
rect 15194 25820 15200 25832
rect 15155 25792 15200 25820
rect 12805 25783 12863 25789
rect 15194 25780 15200 25792
rect 15252 25780 15258 25832
rect 16117 25823 16175 25829
rect 16117 25789 16129 25823
rect 16163 25820 16175 25823
rect 16666 25820 16672 25832
rect 16163 25792 16672 25820
rect 16163 25789 16175 25792
rect 16117 25783 16175 25789
rect 16666 25780 16672 25792
rect 16724 25780 16730 25832
rect 17313 25823 17371 25829
rect 17313 25789 17325 25823
rect 17359 25820 17371 25823
rect 17402 25820 17408 25832
rect 17359 25792 17408 25820
rect 17359 25789 17371 25792
rect 17313 25783 17371 25789
rect 17402 25780 17408 25792
rect 17460 25780 17466 25832
rect 17494 25780 17500 25832
rect 17552 25820 17558 25832
rect 17552 25792 17597 25820
rect 17552 25780 17558 25792
rect 19150 25780 19156 25832
rect 19208 25820 19214 25832
rect 19245 25823 19303 25829
rect 19245 25820 19257 25823
rect 19208 25792 19257 25820
rect 19208 25780 19214 25792
rect 19245 25789 19257 25792
rect 19291 25789 19303 25823
rect 23014 25820 23020 25832
rect 22975 25792 23020 25820
rect 19245 25783 19303 25789
rect 23014 25780 23020 25792
rect 23072 25780 23078 25832
rect 23293 25823 23351 25829
rect 23293 25789 23305 25823
rect 23339 25789 23351 25823
rect 23293 25783 23351 25789
rect 11848 25724 12296 25752
rect 13081 25755 13139 25761
rect 11848 25712 11854 25724
rect 13081 25721 13093 25755
rect 13127 25752 13139 25755
rect 13170 25752 13176 25764
rect 13127 25724 13176 25752
rect 13127 25721 13139 25724
rect 13081 25715 13139 25721
rect 13170 25712 13176 25724
rect 13228 25712 13234 25764
rect 14550 25752 14556 25764
rect 14306 25724 14556 25752
rect 14550 25712 14556 25724
rect 14608 25752 14614 25764
rect 15470 25752 15476 25764
rect 14608 25724 15476 25752
rect 14608 25712 14614 25724
rect 15470 25712 15476 25724
rect 15528 25712 15534 25764
rect 20162 25712 20168 25764
rect 20220 25712 20226 25764
rect 23308 25752 23336 25783
rect 23474 25780 23480 25832
rect 23532 25820 23538 25832
rect 24213 25823 24271 25829
rect 24213 25820 24225 25823
rect 23532 25792 24225 25820
rect 23532 25780 23538 25792
rect 24213 25789 24225 25792
rect 24259 25820 24271 25823
rect 24305 25823 24363 25829
rect 24305 25820 24317 25823
rect 24259 25792 24317 25820
rect 24259 25789 24271 25792
rect 24213 25783 24271 25789
rect 24305 25789 24317 25792
rect 24351 25789 24363 25823
rect 24305 25783 24363 25789
rect 24581 25823 24639 25829
rect 24581 25789 24593 25823
rect 24627 25820 24639 25823
rect 25240 25820 25268 25860
rect 26326 25848 26332 25860
rect 26384 25848 26390 25900
rect 26510 25888 26516 25900
rect 26471 25860 26516 25888
rect 26510 25848 26516 25860
rect 26568 25848 26574 25900
rect 24627 25792 25268 25820
rect 24627 25789 24639 25792
rect 24581 25783 24639 25789
rect 23842 25752 23848 25764
rect 23308 25724 23848 25752
rect 23842 25712 23848 25724
rect 23900 25712 23906 25764
rect 24118 25712 24124 25764
rect 24176 25752 24182 25764
rect 24596 25752 24624 25783
rect 25314 25780 25320 25832
rect 25372 25820 25378 25832
rect 26237 25823 26295 25829
rect 26237 25820 26249 25823
rect 25372 25792 26249 25820
rect 25372 25780 25378 25792
rect 26237 25789 26249 25792
rect 26283 25789 26295 25823
rect 26237 25783 26295 25789
rect 24176 25724 24624 25752
rect 24673 25755 24731 25761
rect 24176 25712 24182 25724
rect 24673 25721 24685 25755
rect 24719 25752 24731 25755
rect 24946 25752 24952 25764
rect 24719 25724 24952 25752
rect 24719 25721 24731 25724
rect 24673 25715 24731 25721
rect 24946 25712 24952 25724
rect 25004 25752 25010 25764
rect 25958 25752 25964 25764
rect 25004 25724 25964 25752
rect 25004 25712 25010 25724
rect 25958 25712 25964 25724
rect 26016 25712 26022 25764
rect 7466 25684 7472 25696
rect 5460 25656 7472 25684
rect 5261 25647 5319 25653
rect 7466 25644 7472 25656
rect 7524 25644 7530 25696
rect 9030 25684 9036 25696
rect 8991 25656 9036 25684
rect 9030 25644 9036 25656
rect 9088 25644 9094 25696
rect 9490 25684 9496 25696
rect 9451 25656 9496 25684
rect 9490 25644 9496 25656
rect 9548 25644 9554 25696
rect 11882 25644 11888 25696
rect 11940 25684 11946 25696
rect 12894 25684 12900 25696
rect 11940 25656 12900 25684
rect 11940 25644 11946 25656
rect 12894 25644 12900 25656
rect 12952 25684 12958 25696
rect 15197 25687 15255 25693
rect 15197 25684 15209 25687
rect 12952 25656 15209 25684
rect 12952 25644 12958 25656
rect 15197 25653 15209 25656
rect 15243 25653 15255 25687
rect 16022 25684 16028 25696
rect 15983 25656 16028 25684
rect 15197 25647 15255 25653
rect 16022 25644 16028 25656
rect 16080 25644 16086 25696
rect 16574 25644 16580 25696
rect 16632 25684 16638 25696
rect 17405 25687 17463 25693
rect 17405 25684 17417 25687
rect 16632 25656 17417 25684
rect 16632 25644 16638 25656
rect 17405 25653 17417 25656
rect 17451 25653 17463 25687
rect 17405 25647 17463 25653
rect 23201 25687 23259 25693
rect 23201 25653 23213 25687
rect 23247 25684 23259 25687
rect 23934 25684 23940 25696
rect 23247 25656 23940 25684
rect 23247 25653 23259 25656
rect 23201 25647 23259 25653
rect 23934 25644 23940 25656
rect 23992 25644 23998 25696
rect 24213 25687 24271 25693
rect 24213 25653 24225 25687
rect 24259 25684 24271 25687
rect 25225 25687 25283 25693
rect 25225 25684 25237 25687
rect 24259 25656 25237 25684
rect 24259 25653 24271 25656
rect 24213 25647 24271 25653
rect 25225 25653 25237 25656
rect 25271 25653 25283 25687
rect 25866 25684 25872 25696
rect 25827 25656 25872 25684
rect 25225 25647 25283 25653
rect 25866 25644 25872 25656
rect 25924 25644 25930 25696
rect 26896 25684 26924 25928
rect 30926 25916 30932 25928
rect 30984 25916 30990 25968
rect 28442 25848 28448 25900
rect 28500 25888 28506 25900
rect 30193 25891 30251 25897
rect 30193 25888 30205 25891
rect 28500 25860 30205 25888
rect 28500 25848 28506 25860
rect 30193 25857 30205 25860
rect 30239 25857 30251 25891
rect 30193 25851 30251 25857
rect 32033 25891 32091 25897
rect 32033 25857 32045 25891
rect 32079 25888 32091 25891
rect 33321 25891 33379 25897
rect 33321 25888 33333 25891
rect 32079 25860 33333 25888
rect 32079 25857 32091 25860
rect 32033 25851 32091 25857
rect 33321 25857 33333 25860
rect 33367 25857 33379 25891
rect 33321 25851 33379 25857
rect 26970 25780 26976 25832
rect 27028 25820 27034 25832
rect 28169 25823 28227 25829
rect 28169 25820 28181 25823
rect 27028 25792 28181 25820
rect 27028 25780 27034 25792
rect 28169 25789 28181 25792
rect 28215 25789 28227 25823
rect 30742 25820 30748 25832
rect 30655 25792 30748 25820
rect 28169 25783 28227 25789
rect 30742 25780 30748 25792
rect 30800 25820 30806 25832
rect 31294 25820 31300 25832
rect 30800 25792 31300 25820
rect 30800 25780 30806 25792
rect 31294 25780 31300 25792
rect 31352 25780 31358 25832
rect 31386 25780 31392 25832
rect 31444 25820 31450 25832
rect 33042 25820 33048 25832
rect 31444 25792 31489 25820
rect 33003 25792 33048 25820
rect 31444 25780 31450 25792
rect 33042 25780 33048 25792
rect 33100 25780 33106 25832
rect 33229 25823 33287 25829
rect 33229 25789 33241 25823
rect 33275 25820 33287 25823
rect 33502 25820 33508 25832
rect 33275 25792 33508 25820
rect 33275 25789 33287 25792
rect 33229 25783 33287 25789
rect 33502 25780 33508 25792
rect 33560 25780 33566 25832
rect 28445 25755 28503 25761
rect 28445 25721 28457 25755
rect 28491 25752 28503 25755
rect 28534 25752 28540 25764
rect 28491 25724 28540 25752
rect 28491 25721 28503 25724
rect 28445 25715 28503 25721
rect 28534 25712 28540 25724
rect 28592 25712 28598 25764
rect 29822 25752 29828 25764
rect 29670 25724 29828 25752
rect 29822 25712 29828 25724
rect 29880 25712 29886 25764
rect 31662 25684 31668 25696
rect 26896 25656 31668 25684
rect 31662 25644 31668 25656
rect 31720 25644 31726 25696
rect 1104 25594 34316 25616
rect 1104 25542 12052 25594
rect 12104 25542 12116 25594
rect 12168 25542 12180 25594
rect 12232 25542 12244 25594
rect 12296 25542 23123 25594
rect 23175 25542 23187 25594
rect 23239 25542 23251 25594
rect 23303 25542 23315 25594
rect 23367 25542 34316 25594
rect 1104 25520 34316 25542
rect 5258 25480 5264 25492
rect 4724 25452 5264 25480
rect 2958 25412 2964 25424
rect 1964 25384 2964 25412
rect 1762 25344 1768 25356
rect 1723 25316 1768 25344
rect 1762 25304 1768 25316
rect 1820 25304 1826 25356
rect 1964 25353 1992 25384
rect 2958 25372 2964 25384
rect 3016 25372 3022 25424
rect 1949 25347 2007 25353
rect 1949 25313 1961 25347
rect 1995 25313 2007 25347
rect 2501 25347 2559 25353
rect 2501 25344 2513 25347
rect 1949 25307 2007 25313
rect 2240 25316 2513 25344
rect 1857 25279 1915 25285
rect 1857 25245 1869 25279
rect 1903 25276 1915 25279
rect 2240 25276 2268 25316
rect 2501 25313 2513 25316
rect 2547 25313 2559 25347
rect 2501 25307 2559 25313
rect 2593 25347 2651 25353
rect 2593 25313 2605 25347
rect 2639 25344 2651 25347
rect 3326 25344 3332 25356
rect 2639 25316 3332 25344
rect 2639 25313 2651 25316
rect 2593 25307 2651 25313
rect 3326 25304 3332 25316
rect 3384 25304 3390 25356
rect 4724 25353 4752 25452
rect 5258 25440 5264 25452
rect 5316 25440 5322 25492
rect 8113 25483 8171 25489
rect 8113 25449 8125 25483
rect 8159 25480 8171 25483
rect 8294 25480 8300 25492
rect 8159 25452 8300 25480
rect 8159 25449 8171 25452
rect 8113 25443 8171 25449
rect 8294 25440 8300 25452
rect 8352 25480 8358 25492
rect 12618 25480 12624 25492
rect 8352 25452 12624 25480
rect 8352 25440 8358 25452
rect 12618 25440 12624 25452
rect 12676 25440 12682 25492
rect 13081 25483 13139 25489
rect 13081 25449 13093 25483
rect 13127 25480 13139 25483
rect 13170 25480 13176 25492
rect 13127 25452 13176 25480
rect 13127 25449 13139 25452
rect 13081 25443 13139 25449
rect 13170 25440 13176 25452
rect 13228 25440 13234 25492
rect 15105 25483 15163 25489
rect 15105 25449 15117 25483
rect 15151 25480 15163 25483
rect 25314 25480 25320 25492
rect 15151 25452 24256 25480
rect 15151 25449 15163 25452
rect 15105 25443 15163 25449
rect 5031 25415 5089 25421
rect 5031 25381 5043 25415
rect 5077 25412 5089 25415
rect 5534 25412 5540 25424
rect 5077 25384 5540 25412
rect 5077 25381 5089 25384
rect 5031 25375 5089 25381
rect 5534 25372 5540 25384
rect 5592 25372 5598 25424
rect 7006 25412 7012 25424
rect 6670 25384 7012 25412
rect 7006 25372 7012 25384
rect 7064 25372 7070 25424
rect 9490 25372 9496 25424
rect 9548 25412 9554 25424
rect 9677 25415 9735 25421
rect 9677 25412 9689 25415
rect 9548 25384 9689 25412
rect 9548 25372 9554 25384
rect 9677 25381 9689 25384
rect 9723 25381 9735 25415
rect 9677 25375 9735 25381
rect 12802 25372 12808 25424
rect 12860 25412 12866 25424
rect 12860 25384 12905 25412
rect 12860 25372 12866 25384
rect 18782 25372 18788 25424
rect 18840 25412 18846 25424
rect 23934 25412 23940 25424
rect 18840 25384 23796 25412
rect 23895 25384 23940 25412
rect 18840 25372 18846 25384
rect 4709 25347 4767 25353
rect 4709 25313 4721 25347
rect 4755 25313 4767 25347
rect 4709 25307 4767 25313
rect 4801 25347 4859 25353
rect 4801 25313 4813 25347
rect 4847 25313 4859 25347
rect 4801 25307 4859 25313
rect 1903 25248 2268 25276
rect 2685 25279 2743 25285
rect 1903 25245 1915 25248
rect 1857 25239 1915 25245
rect 2685 25245 2697 25279
rect 2731 25245 2743 25279
rect 2685 25239 2743 25245
rect 2700 25208 2728 25239
rect 2774 25236 2780 25288
rect 2832 25276 2838 25288
rect 2832 25248 2877 25276
rect 2832 25236 2838 25248
rect 2958 25236 2964 25288
rect 3016 25236 3022 25288
rect 2976 25208 3004 25236
rect 2700 25180 3004 25208
rect 4816 25208 4844 25307
rect 4890 25304 4896 25356
rect 4948 25344 4954 25356
rect 4948 25316 4993 25344
rect 4948 25304 4954 25316
rect 7374 25304 7380 25356
rect 7432 25344 7438 25356
rect 7926 25344 7932 25356
rect 7432 25316 7477 25344
rect 7887 25316 7932 25344
rect 7432 25304 7438 25316
rect 7926 25304 7932 25316
rect 7984 25304 7990 25356
rect 9858 25344 9864 25356
rect 9819 25316 9864 25344
rect 9858 25304 9864 25316
rect 9916 25304 9922 25356
rect 10870 25344 10876 25356
rect 10831 25316 10876 25344
rect 10870 25304 10876 25316
rect 10928 25304 10934 25356
rect 11146 25344 11152 25356
rect 11107 25316 11152 25344
rect 11146 25304 11152 25316
rect 11204 25304 11210 25356
rect 11241 25347 11299 25353
rect 11241 25313 11253 25347
rect 11287 25344 11299 25347
rect 11422 25344 11428 25356
rect 11287 25316 11428 25344
rect 11287 25313 11299 25316
rect 11241 25307 11299 25313
rect 11422 25304 11428 25316
rect 11480 25304 11486 25356
rect 12434 25344 12440 25356
rect 12395 25316 12440 25344
rect 12434 25304 12440 25316
rect 12492 25304 12498 25356
rect 12526 25304 12532 25356
rect 12584 25344 12590 25356
rect 12713 25347 12771 25353
rect 12584 25316 12629 25344
rect 12584 25304 12590 25316
rect 12713 25313 12725 25347
rect 12759 25313 12771 25347
rect 12713 25307 12771 25313
rect 5166 25276 5172 25288
rect 5127 25248 5172 25276
rect 5166 25236 5172 25248
rect 5224 25236 5230 25288
rect 7098 25276 7104 25288
rect 7059 25248 7104 25276
rect 7098 25236 7104 25248
rect 7156 25236 7162 25288
rect 4816 25180 5672 25208
rect 5644 25152 5672 25180
rect 7466 25168 7472 25220
rect 7524 25208 7530 25220
rect 7524 25180 9628 25208
rect 7524 25168 7530 25180
rect 2958 25140 2964 25152
rect 2919 25112 2964 25140
rect 2958 25100 2964 25112
rect 3016 25100 3022 25152
rect 4430 25100 4436 25152
rect 4488 25140 4494 25152
rect 4525 25143 4583 25149
rect 4525 25140 4537 25143
rect 4488 25112 4537 25140
rect 4488 25100 4494 25112
rect 4525 25109 4537 25112
rect 4571 25109 4583 25143
rect 5626 25140 5632 25152
rect 5587 25112 5632 25140
rect 4525 25103 4583 25109
rect 5626 25100 5632 25112
rect 5684 25100 5690 25152
rect 9490 25140 9496 25152
rect 9451 25112 9496 25140
rect 9490 25100 9496 25112
rect 9548 25100 9554 25152
rect 9600 25140 9628 25180
rect 10042 25168 10048 25220
rect 10100 25208 10106 25220
rect 10597 25211 10655 25217
rect 10597 25208 10609 25211
rect 10100 25180 10609 25208
rect 10100 25168 10106 25180
rect 10597 25177 10609 25180
rect 10643 25177 10655 25211
rect 10597 25171 10655 25177
rect 12158 25168 12164 25220
rect 12216 25208 12222 25220
rect 12728 25208 12756 25307
rect 12894 25304 12900 25356
rect 12952 25344 12958 25356
rect 15464 25347 15522 25353
rect 12952 25316 12997 25344
rect 12952 25304 12958 25316
rect 15464 25313 15476 25347
rect 15510 25344 15522 25347
rect 16206 25344 16212 25356
rect 15510 25316 16212 25344
rect 15510 25313 15522 25316
rect 15464 25307 15522 25313
rect 16206 25304 16212 25316
rect 16264 25304 16270 25356
rect 18138 25304 18144 25356
rect 18196 25344 18202 25356
rect 18702 25347 18760 25353
rect 18702 25344 18714 25347
rect 18196 25316 18714 25344
rect 18196 25304 18202 25316
rect 18702 25313 18714 25316
rect 18748 25313 18760 25347
rect 18702 25307 18760 25313
rect 22922 25304 22928 25356
rect 22980 25344 22986 25356
rect 23201 25347 23259 25353
rect 23201 25344 23213 25347
rect 22980 25316 23213 25344
rect 22980 25304 22986 25316
rect 23201 25313 23213 25316
rect 23247 25313 23259 25347
rect 23474 25344 23480 25356
rect 23435 25316 23480 25344
rect 23201 25307 23259 25313
rect 23474 25304 23480 25316
rect 23532 25304 23538 25356
rect 23768 25344 23796 25384
rect 23934 25372 23940 25384
rect 23992 25372 23998 25424
rect 24118 25344 24124 25356
rect 23768 25316 24124 25344
rect 24118 25304 24124 25316
rect 24176 25304 24182 25356
rect 13814 25236 13820 25288
rect 13872 25276 13878 25288
rect 14918 25276 14924 25288
rect 13872 25248 14924 25276
rect 13872 25236 13878 25248
rect 14918 25236 14924 25248
rect 14976 25276 14982 25288
rect 15197 25279 15255 25285
rect 15197 25276 15209 25279
rect 14976 25248 15209 25276
rect 14976 25236 14982 25248
rect 15197 25245 15209 25248
rect 15243 25245 15255 25279
rect 15197 25239 15255 25245
rect 18969 25279 19027 25285
rect 18969 25245 18981 25279
rect 19015 25276 19027 25279
rect 19150 25276 19156 25288
rect 19015 25248 19156 25276
rect 19015 25245 19027 25248
rect 18969 25239 19027 25245
rect 19150 25236 19156 25248
rect 19208 25236 19214 25288
rect 13722 25208 13728 25220
rect 12216 25180 13728 25208
rect 12216 25168 12222 25180
rect 13722 25168 13728 25180
rect 13780 25168 13786 25220
rect 17494 25168 17500 25220
rect 17552 25168 17558 25220
rect 15105 25143 15163 25149
rect 15105 25140 15117 25143
rect 9600 25112 15117 25140
rect 15105 25109 15117 25112
rect 15151 25109 15163 25143
rect 15105 25103 15163 25109
rect 16577 25143 16635 25149
rect 16577 25109 16589 25143
rect 16623 25140 16635 25143
rect 16666 25140 16672 25152
rect 16623 25112 16672 25140
rect 16623 25109 16635 25112
rect 16577 25103 16635 25109
rect 16666 25100 16672 25112
rect 16724 25100 16730 25152
rect 17126 25100 17132 25152
rect 17184 25140 17190 25152
rect 17512 25140 17540 25168
rect 17589 25143 17647 25149
rect 17589 25140 17601 25143
rect 17184 25112 17601 25140
rect 17184 25100 17190 25112
rect 17589 25109 17601 25112
rect 17635 25109 17647 25143
rect 17589 25103 17647 25109
rect 23385 25143 23443 25149
rect 23385 25109 23397 25143
rect 23431 25140 23443 25143
rect 23842 25140 23848 25152
rect 23431 25112 23848 25140
rect 23431 25109 23443 25112
rect 23385 25103 23443 25109
rect 23842 25100 23848 25112
rect 23900 25100 23906 25152
rect 24228 25140 24256 25452
rect 24320 25452 25320 25480
rect 24320 25353 24348 25452
rect 25314 25440 25320 25452
rect 25372 25480 25378 25492
rect 25409 25483 25467 25489
rect 25409 25480 25421 25483
rect 25372 25452 25421 25480
rect 25372 25440 25378 25452
rect 25409 25449 25421 25452
rect 25455 25449 25467 25483
rect 28534 25480 28540 25492
rect 28495 25452 28540 25480
rect 25409 25443 25467 25449
rect 28534 25440 28540 25452
rect 28592 25440 28598 25492
rect 29457 25483 29515 25489
rect 29457 25449 29469 25483
rect 29503 25480 29515 25483
rect 31386 25480 31392 25492
rect 29503 25452 31392 25480
rect 29503 25449 29515 25452
rect 29457 25443 29515 25449
rect 31386 25440 31392 25452
rect 31444 25440 31450 25492
rect 25866 25372 25872 25424
rect 25924 25412 25930 25424
rect 26522 25415 26580 25421
rect 26522 25412 26534 25415
rect 25924 25384 26534 25412
rect 25924 25372 25930 25384
rect 26522 25381 26534 25384
rect 26568 25381 26580 25415
rect 26522 25375 26580 25381
rect 29564 25384 31616 25412
rect 24305 25347 24363 25353
rect 24305 25313 24317 25347
rect 24351 25313 24363 25347
rect 28166 25344 28172 25356
rect 28127 25316 28172 25344
rect 24305 25307 24363 25313
rect 28166 25304 28172 25316
rect 28224 25304 28230 25356
rect 28323 25347 28381 25353
rect 28323 25313 28335 25347
rect 28369 25344 28381 25347
rect 28442 25344 28448 25356
rect 28369 25316 28448 25344
rect 28369 25313 28381 25316
rect 28323 25307 28381 25313
rect 28442 25304 28448 25316
rect 28500 25304 28506 25356
rect 29362 25344 29368 25356
rect 29275 25316 29368 25344
rect 29362 25304 29368 25316
rect 29420 25304 29426 25356
rect 29564 25353 29592 25384
rect 31588 25356 31616 25384
rect 31662 25372 31668 25424
rect 31720 25412 31726 25424
rect 32953 25415 33011 25421
rect 32953 25412 32965 25415
rect 31720 25384 32965 25412
rect 31720 25372 31726 25384
rect 32953 25381 32965 25384
rect 32999 25381 33011 25415
rect 32953 25375 33011 25381
rect 29549 25347 29607 25353
rect 29549 25313 29561 25347
rect 29595 25313 29607 25347
rect 29549 25307 29607 25313
rect 30929 25347 30987 25353
rect 30929 25313 30941 25347
rect 30975 25313 30987 25347
rect 31570 25344 31576 25356
rect 31531 25316 31576 25344
rect 30929 25307 30987 25313
rect 26789 25279 26847 25285
rect 26789 25245 26801 25279
rect 26835 25276 26847 25279
rect 26878 25276 26884 25288
rect 26835 25248 26884 25276
rect 26835 25245 26847 25248
rect 26789 25239 26847 25245
rect 26878 25236 26884 25248
rect 26936 25236 26942 25288
rect 29380 25276 29408 25304
rect 30944 25276 30972 25307
rect 31570 25304 31576 25316
rect 31628 25304 31634 25356
rect 31754 25344 31760 25356
rect 31715 25316 31760 25344
rect 31754 25304 31760 25316
rect 31812 25304 31818 25356
rect 32217 25347 32275 25353
rect 32217 25313 32229 25347
rect 32263 25344 32275 25347
rect 33318 25344 33324 25356
rect 32263 25316 33324 25344
rect 32263 25313 32275 25316
rect 32217 25307 32275 25313
rect 33318 25304 33324 25316
rect 33376 25304 33382 25356
rect 33502 25344 33508 25356
rect 33463 25316 33508 25344
rect 33502 25304 33508 25316
rect 33560 25304 33566 25356
rect 29380 25248 30972 25276
rect 31846 25168 31852 25220
rect 31904 25208 31910 25220
rect 32309 25211 32367 25217
rect 32309 25208 32321 25211
rect 31904 25180 32321 25208
rect 31904 25168 31910 25180
rect 32309 25177 32321 25180
rect 32355 25177 32367 25211
rect 32309 25171 32367 25177
rect 33134 25140 33140 25152
rect 24228 25112 33140 25140
rect 33134 25100 33140 25112
rect 33192 25100 33198 25152
rect 1104 25050 34316 25072
rect 1104 24998 6517 25050
rect 6569 24998 6581 25050
rect 6633 24998 6645 25050
rect 6697 24998 6709 25050
rect 6761 24998 17588 25050
rect 17640 24998 17652 25050
rect 17704 24998 17716 25050
rect 17768 24998 17780 25050
rect 17832 24998 28658 25050
rect 28710 24998 28722 25050
rect 28774 24998 28786 25050
rect 28838 24998 28850 25050
rect 28902 24998 34316 25050
rect 1104 24976 34316 24998
rect 4890 24896 4896 24948
rect 4948 24936 4954 24948
rect 5169 24939 5227 24945
rect 5169 24936 5181 24939
rect 4948 24908 5181 24936
rect 4948 24896 4954 24908
rect 5169 24905 5181 24908
rect 5215 24905 5227 24939
rect 5169 24899 5227 24905
rect 6825 24939 6883 24945
rect 6825 24905 6837 24939
rect 6871 24936 6883 24939
rect 7098 24936 7104 24948
rect 6871 24908 7104 24936
rect 6871 24905 6883 24908
rect 6825 24899 6883 24905
rect 7098 24896 7104 24908
rect 7156 24896 7162 24948
rect 7282 24896 7288 24948
rect 7340 24936 7346 24948
rect 8297 24939 8355 24945
rect 8297 24936 8309 24939
rect 7340 24908 8309 24936
rect 7340 24896 7346 24908
rect 8297 24905 8309 24908
rect 8343 24936 8355 24939
rect 8343 24908 9720 24936
rect 8343 24905 8355 24908
rect 8297 24899 8355 24905
rect 9582 24868 9588 24880
rect 7484 24840 9588 24868
rect 5074 24760 5080 24812
rect 5132 24800 5138 24812
rect 5132 24772 5396 24800
rect 5132 24760 5138 24772
rect 1486 24692 1492 24744
rect 1544 24732 1550 24744
rect 2777 24735 2835 24741
rect 2777 24732 2789 24735
rect 1544 24704 2789 24732
rect 1544 24692 1550 24704
rect 2777 24701 2789 24704
rect 2823 24732 2835 24735
rect 2823 24704 3464 24732
rect 2823 24701 2835 24704
rect 2777 24695 2835 24701
rect 2532 24667 2590 24673
rect 2532 24633 2544 24667
rect 2578 24664 2590 24667
rect 2958 24664 2964 24676
rect 2578 24636 2964 24664
rect 2578 24633 2590 24636
rect 2532 24627 2590 24633
rect 2958 24624 2964 24636
rect 3016 24624 3022 24676
rect 3436 24664 3464 24704
rect 4430 24692 4436 24744
rect 4488 24741 4494 24744
rect 5368 24741 5396 24772
rect 5626 24760 5632 24812
rect 5684 24800 5690 24812
rect 7484 24809 7512 24840
rect 9582 24828 9588 24840
rect 9640 24828 9646 24880
rect 9692 24868 9720 24908
rect 9766 24896 9772 24948
rect 9824 24936 9830 24948
rect 10226 24936 10232 24948
rect 9824 24908 10232 24936
rect 9824 24896 9830 24908
rect 10226 24896 10232 24908
rect 10284 24936 10290 24948
rect 15010 24936 15016 24948
rect 10284 24908 15016 24936
rect 10284 24896 10290 24908
rect 15010 24896 15016 24908
rect 15068 24896 15074 24948
rect 16206 24936 16212 24948
rect 16167 24908 16212 24936
rect 16206 24896 16212 24908
rect 16264 24896 16270 24948
rect 30742 24936 30748 24948
rect 30703 24908 30748 24936
rect 30742 24896 30748 24908
rect 30800 24896 30806 24948
rect 12158 24868 12164 24880
rect 9692 24840 12164 24868
rect 7285 24803 7343 24809
rect 7285 24800 7297 24803
rect 5684 24772 7297 24800
rect 5684 24760 5690 24772
rect 7285 24769 7297 24772
rect 7331 24769 7343 24803
rect 7285 24763 7343 24769
rect 7469 24803 7527 24809
rect 7469 24769 7481 24803
rect 7515 24769 7527 24803
rect 7469 24763 7527 24769
rect 9401 24803 9459 24809
rect 9401 24769 9413 24803
rect 9447 24800 9459 24803
rect 9692 24800 9720 24840
rect 12158 24828 12164 24840
rect 12216 24828 12222 24880
rect 13998 24828 14004 24880
rect 14056 24868 14062 24880
rect 14918 24868 14924 24880
rect 14056 24840 14924 24868
rect 14056 24828 14062 24840
rect 14918 24828 14924 24840
rect 14976 24828 14982 24880
rect 10778 24800 10784 24812
rect 9447 24772 9720 24800
rect 10739 24772 10784 24800
rect 9447 24769 9459 24772
rect 9401 24763 9459 24769
rect 10778 24760 10784 24772
rect 10836 24760 10842 24812
rect 11882 24760 11888 24812
rect 11940 24800 11946 24812
rect 12069 24803 12127 24809
rect 12069 24800 12081 24803
rect 11940 24772 12081 24800
rect 11940 24760 11946 24772
rect 12069 24769 12081 24772
rect 12115 24769 12127 24803
rect 12069 24763 12127 24769
rect 15565 24803 15623 24809
rect 15565 24769 15577 24803
rect 15611 24800 15623 24803
rect 16298 24800 16304 24812
rect 15611 24772 16160 24800
rect 16259 24772 16304 24800
rect 15611 24769 15623 24772
rect 15565 24763 15623 24769
rect 4488 24732 4500 24741
rect 4709 24735 4767 24741
rect 4488 24704 4533 24732
rect 4488 24695 4500 24704
rect 4709 24701 4721 24735
rect 4755 24701 4767 24735
rect 5169 24735 5227 24741
rect 5169 24732 5181 24735
rect 4709 24695 4767 24701
rect 5092 24704 5181 24732
rect 4488 24692 4494 24695
rect 4724 24664 4752 24695
rect 5092 24676 5120 24704
rect 5169 24701 5181 24704
rect 5215 24701 5227 24735
rect 5169 24695 5227 24701
rect 5353 24735 5411 24741
rect 5353 24701 5365 24735
rect 5399 24701 5411 24735
rect 7190 24732 7196 24744
rect 7151 24704 7196 24732
rect 5353 24695 5411 24701
rect 7190 24692 7196 24704
rect 7248 24692 7254 24744
rect 8294 24732 8300 24744
rect 8255 24704 8300 24732
rect 8294 24692 8300 24704
rect 8352 24692 8358 24744
rect 9217 24735 9275 24741
rect 9217 24701 9229 24735
rect 9263 24732 9275 24735
rect 9490 24732 9496 24744
rect 9263 24704 9496 24732
rect 9263 24701 9275 24704
rect 9217 24695 9275 24701
rect 9490 24692 9496 24704
rect 9548 24692 9554 24744
rect 10226 24732 10232 24744
rect 10187 24704 10232 24732
rect 10226 24692 10232 24704
rect 10284 24692 10290 24744
rect 10689 24735 10747 24741
rect 10689 24701 10701 24735
rect 10735 24701 10747 24735
rect 10689 24695 10747 24701
rect 10873 24735 10931 24741
rect 10873 24701 10885 24735
rect 10919 24701 10931 24735
rect 12250 24732 12256 24744
rect 12211 24704 12256 24732
rect 10873 24695 10931 24701
rect 3436 24636 4752 24664
rect 5074 24624 5080 24676
rect 5132 24624 5138 24676
rect 9309 24667 9367 24673
rect 9309 24633 9321 24667
rect 9355 24664 9367 24667
rect 9398 24664 9404 24676
rect 9355 24636 9404 24664
rect 9355 24633 9367 24636
rect 9309 24627 9367 24633
rect 9398 24624 9404 24636
rect 9456 24624 9462 24676
rect 9950 24624 9956 24676
rect 10008 24664 10014 24676
rect 10704 24664 10732 24695
rect 10008 24636 10732 24664
rect 10888 24664 10916 24695
rect 12250 24692 12256 24704
rect 12308 24692 12314 24744
rect 12345 24735 12403 24741
rect 12345 24701 12357 24735
rect 12391 24732 12403 24735
rect 12986 24732 12992 24744
rect 12391 24704 12992 24732
rect 12391 24701 12403 24704
rect 12345 24695 12403 24701
rect 12986 24692 12992 24704
rect 13044 24692 13050 24744
rect 13630 24732 13636 24744
rect 13591 24704 13636 24732
rect 13630 24692 13636 24704
rect 13688 24692 13694 24744
rect 15286 24732 15292 24744
rect 15247 24704 15292 24732
rect 15286 24692 15292 24704
rect 15344 24692 15350 24744
rect 16022 24732 16028 24744
rect 15983 24704 16028 24732
rect 16022 24692 16028 24704
rect 16080 24692 16086 24744
rect 16132 24741 16160 24772
rect 16298 24760 16304 24772
rect 16356 24760 16362 24812
rect 16666 24760 16672 24812
rect 16724 24800 16730 24812
rect 18877 24803 18935 24809
rect 16724 24772 18000 24800
rect 16724 24760 16730 24772
rect 16117 24735 16175 24741
rect 16117 24701 16129 24735
rect 16163 24732 16175 24735
rect 16574 24732 16580 24744
rect 16163 24704 16580 24732
rect 16163 24701 16175 24704
rect 16117 24695 16175 24701
rect 16574 24692 16580 24704
rect 16632 24692 16638 24744
rect 17402 24692 17408 24744
rect 17460 24732 17466 24744
rect 17972 24741 18000 24772
rect 18877 24769 18889 24803
rect 18923 24800 18935 24803
rect 19150 24800 19156 24812
rect 18923 24772 19156 24800
rect 18923 24769 18935 24772
rect 18877 24763 18935 24769
rect 19150 24760 19156 24772
rect 19208 24800 19214 24812
rect 20162 24800 20168 24812
rect 19208 24772 20168 24800
rect 19208 24760 19214 24772
rect 20162 24760 20168 24772
rect 20220 24760 20226 24812
rect 22922 24800 22928 24812
rect 21284 24772 22928 24800
rect 17497 24735 17555 24741
rect 17497 24732 17509 24735
rect 17460 24704 17509 24732
rect 17460 24692 17466 24704
rect 17497 24701 17509 24704
rect 17543 24701 17555 24735
rect 17497 24695 17555 24701
rect 17773 24735 17831 24741
rect 17773 24701 17785 24735
rect 17819 24701 17831 24735
rect 17773 24695 17831 24701
rect 17957 24735 18015 24741
rect 17957 24701 17969 24735
rect 18003 24701 18015 24735
rect 21082 24732 21088 24744
rect 17957 24695 18015 24701
rect 20364 24704 21088 24732
rect 13354 24664 13360 24676
rect 10888 24636 13360 24664
rect 10008 24624 10014 24636
rect 13354 24624 13360 24636
rect 13412 24624 13418 24676
rect 14366 24624 14372 24676
rect 14424 24664 14430 24676
rect 14829 24667 14887 24673
rect 14829 24664 14841 24667
rect 14424 24636 14841 24664
rect 14424 24624 14430 24636
rect 14829 24633 14841 24636
rect 14875 24664 14887 24667
rect 15194 24664 15200 24676
rect 14875 24636 15200 24664
rect 14875 24633 14887 24636
rect 14829 24627 14887 24633
rect 15194 24624 15200 24636
rect 15252 24624 15258 24676
rect 15381 24667 15439 24673
rect 15381 24633 15393 24667
rect 15427 24664 15439 24667
rect 16040 24664 16068 24692
rect 15427 24636 16068 24664
rect 15427 24633 15439 24636
rect 15381 24627 15439 24633
rect 17126 24624 17132 24676
rect 17184 24664 17190 24676
rect 17788 24664 17816 24695
rect 17184 24636 17816 24664
rect 19153 24667 19211 24673
rect 17184 24624 17190 24636
rect 19153 24633 19165 24667
rect 19199 24664 19211 24667
rect 19426 24664 19432 24676
rect 19199 24636 19432 24664
rect 19199 24633 19211 24636
rect 19153 24627 19211 24633
rect 19426 24624 19432 24636
rect 19484 24624 19490 24676
rect 1397 24599 1455 24605
rect 1397 24565 1409 24599
rect 1443 24596 1455 24599
rect 2130 24596 2136 24608
rect 1443 24568 2136 24596
rect 1443 24565 1455 24568
rect 1397 24559 1455 24565
rect 2130 24556 2136 24568
rect 2188 24556 2194 24608
rect 3326 24596 3332 24608
rect 3239 24568 3332 24596
rect 3326 24556 3332 24568
rect 3384 24596 3390 24608
rect 5166 24596 5172 24608
rect 3384 24568 5172 24596
rect 3384 24556 3390 24568
rect 5166 24556 5172 24568
rect 5224 24556 5230 24608
rect 8846 24596 8852 24608
rect 8807 24568 8852 24596
rect 8846 24556 8852 24568
rect 8904 24556 8910 24608
rect 9858 24556 9864 24608
rect 9916 24596 9922 24608
rect 10137 24599 10195 24605
rect 10137 24596 10149 24599
rect 9916 24568 10149 24596
rect 9916 24556 9922 24568
rect 10137 24565 10149 24568
rect 10183 24565 10195 24599
rect 10137 24559 10195 24565
rect 11238 24556 11244 24608
rect 11296 24596 11302 24608
rect 12069 24599 12127 24605
rect 12069 24596 12081 24599
rect 11296 24568 12081 24596
rect 11296 24556 11302 24568
rect 12069 24565 12081 24568
rect 12115 24565 12127 24599
rect 13814 24596 13820 24608
rect 13775 24568 13820 24596
rect 12069 24559 12127 24565
rect 13814 24556 13820 24568
rect 13872 24556 13878 24608
rect 17218 24556 17224 24608
rect 17276 24596 17282 24608
rect 17313 24599 17371 24605
rect 17313 24596 17325 24599
rect 17276 24568 17325 24596
rect 17276 24556 17282 24568
rect 17313 24565 17325 24568
rect 17359 24565 17371 24599
rect 17313 24559 17371 24565
rect 19518 24556 19524 24608
rect 19576 24596 19582 24608
rect 20364 24596 20392 24704
rect 21082 24692 21088 24704
rect 21140 24692 21146 24744
rect 21284 24741 21312 24772
rect 22922 24760 22928 24772
rect 22980 24760 22986 24812
rect 23474 24800 23480 24812
rect 23435 24772 23480 24800
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 30466 24800 30472 24812
rect 29932 24772 30472 24800
rect 21269 24735 21327 24741
rect 21269 24701 21281 24735
rect 21315 24701 21327 24735
rect 21269 24695 21327 24701
rect 21545 24735 21603 24741
rect 21545 24701 21557 24735
rect 21591 24732 21603 24735
rect 22649 24735 22707 24741
rect 21591 24704 22094 24732
rect 21591 24701 21603 24704
rect 21545 24695 21603 24701
rect 20438 24624 20444 24676
rect 20496 24664 20502 24676
rect 21453 24667 21511 24673
rect 21453 24664 21465 24667
rect 20496 24636 21465 24664
rect 20496 24624 20502 24636
rect 21453 24633 21465 24636
rect 21499 24633 21511 24667
rect 22066 24664 22094 24704
rect 22649 24701 22661 24735
rect 22695 24732 22707 24735
rect 23569 24735 23627 24741
rect 22695 24704 23520 24732
rect 22695 24701 22707 24704
rect 22649 24695 22707 24701
rect 23014 24664 23020 24676
rect 22066 24636 23020 24664
rect 21453 24627 21511 24633
rect 23014 24624 23020 24636
rect 23072 24624 23078 24676
rect 19576 24568 20392 24596
rect 19576 24556 19582 24568
rect 20530 24556 20536 24608
rect 20588 24596 20594 24608
rect 20625 24599 20683 24605
rect 20625 24596 20637 24599
rect 20588 24568 20637 24596
rect 20588 24556 20594 24568
rect 20625 24565 20637 24568
rect 20671 24565 20683 24599
rect 20625 24559 20683 24565
rect 20806 24556 20812 24608
rect 20864 24596 20870 24608
rect 21361 24599 21419 24605
rect 21361 24596 21373 24599
rect 20864 24568 21373 24596
rect 20864 24556 20870 24568
rect 21361 24565 21373 24568
rect 21407 24565 21419 24599
rect 21361 24559 21419 24565
rect 22554 24556 22560 24608
rect 22612 24596 22618 24608
rect 22741 24599 22799 24605
rect 22741 24596 22753 24599
rect 22612 24568 22753 24596
rect 22612 24556 22618 24568
rect 22741 24565 22753 24568
rect 22787 24565 22799 24599
rect 23492 24596 23520 24704
rect 23569 24701 23581 24735
rect 23615 24701 23627 24735
rect 23750 24732 23756 24744
rect 23711 24704 23756 24732
rect 23569 24695 23627 24701
rect 23584 24664 23612 24695
rect 23750 24692 23756 24704
rect 23808 24692 23814 24744
rect 23934 24692 23940 24744
rect 23992 24732 23998 24744
rect 24121 24735 24179 24741
rect 24121 24732 24133 24735
rect 23992 24704 24133 24732
rect 23992 24692 23998 24704
rect 24121 24701 24133 24704
rect 24167 24701 24179 24735
rect 25038 24732 25044 24744
rect 24999 24704 25044 24732
rect 24121 24695 24179 24701
rect 25038 24692 25044 24704
rect 25096 24692 25102 24744
rect 27985 24735 28043 24741
rect 27985 24701 27997 24735
rect 28031 24732 28043 24735
rect 28166 24732 28172 24744
rect 28031 24704 28172 24732
rect 28031 24701 28043 24704
rect 27985 24695 28043 24701
rect 28166 24692 28172 24704
rect 28224 24692 28230 24744
rect 28261 24735 28319 24741
rect 28261 24701 28273 24735
rect 28307 24732 28319 24735
rect 29178 24732 29184 24744
rect 28307 24704 29184 24732
rect 28307 24701 28319 24704
rect 28261 24695 28319 24701
rect 29178 24692 29184 24704
rect 29236 24692 29242 24744
rect 29932 24741 29960 24772
rect 30466 24760 30472 24772
rect 30524 24800 30530 24812
rect 30926 24800 30932 24812
rect 30524 24772 30932 24800
rect 30524 24760 30530 24772
rect 30926 24760 30932 24772
rect 30984 24760 30990 24812
rect 33318 24800 33324 24812
rect 33279 24772 33324 24800
rect 33318 24760 33324 24772
rect 33376 24760 33382 24812
rect 29733 24735 29791 24741
rect 29733 24701 29745 24735
rect 29779 24701 29791 24735
rect 29733 24695 29791 24701
rect 29917 24735 29975 24741
rect 29917 24701 29929 24735
rect 29963 24701 29975 24735
rect 29917 24695 29975 24701
rect 30285 24735 30343 24741
rect 30285 24701 30297 24735
rect 30331 24732 30343 24735
rect 30742 24732 30748 24744
rect 30331 24704 30748 24732
rect 30331 24701 30343 24704
rect 30285 24695 30343 24701
rect 23842 24664 23848 24676
rect 23584 24636 23848 24664
rect 23842 24624 23848 24636
rect 23900 24624 23906 24676
rect 26418 24664 26424 24676
rect 23952 24636 26424 24664
rect 23952 24596 23980 24636
rect 26418 24624 26424 24636
rect 26476 24624 26482 24676
rect 29748 24664 29776 24695
rect 30742 24692 30748 24704
rect 30800 24692 30806 24744
rect 32122 24732 32128 24744
rect 32083 24704 32128 24732
rect 32122 24692 32128 24704
rect 32180 24692 32186 24744
rect 32950 24692 32956 24744
rect 33008 24732 33014 24744
rect 33045 24735 33103 24741
rect 33045 24732 33057 24735
rect 33008 24704 33057 24732
rect 33008 24692 33014 24704
rect 33045 24701 33057 24704
rect 33091 24701 33103 24735
rect 33226 24732 33232 24744
rect 33187 24704 33232 24732
rect 33045 24695 33103 24701
rect 33226 24692 33232 24704
rect 33284 24692 33290 24744
rect 31754 24664 31760 24676
rect 29748 24636 31760 24664
rect 31754 24624 31760 24636
rect 31812 24624 31818 24676
rect 31880 24667 31938 24673
rect 31880 24633 31892 24667
rect 31926 24664 31938 24667
rect 32968 24664 32996 24692
rect 31926 24636 32996 24664
rect 31926 24633 31938 24636
rect 31880 24627 31938 24633
rect 25222 24596 25228 24608
rect 23492 24568 23980 24596
rect 25183 24568 25228 24596
rect 22741 24559 22799 24565
rect 25222 24556 25228 24568
rect 25280 24556 25286 24608
rect 27154 24556 27160 24608
rect 27212 24596 27218 24608
rect 28083 24599 28141 24605
rect 28083 24596 28095 24599
rect 27212 24568 28095 24596
rect 27212 24556 27218 24568
rect 28083 24565 28095 24568
rect 28129 24565 28141 24599
rect 28083 24559 28141 24565
rect 28169 24599 28227 24605
rect 28169 24565 28181 24599
rect 28215 24596 28227 24599
rect 28258 24596 28264 24608
rect 28215 24568 28264 24596
rect 28215 24565 28227 24568
rect 28169 24559 28227 24565
rect 28258 24556 28264 24568
rect 28316 24556 28322 24608
rect 28350 24556 28356 24608
rect 28408 24596 28414 24608
rect 29917 24599 29975 24605
rect 29917 24596 29929 24599
rect 28408 24568 29929 24596
rect 28408 24556 28414 24568
rect 29917 24565 29929 24568
rect 29963 24565 29975 24599
rect 29917 24559 29975 24565
rect 1104 24506 34316 24528
rect 1104 24454 12052 24506
rect 12104 24454 12116 24506
rect 12168 24454 12180 24506
rect 12232 24454 12244 24506
rect 12296 24454 23123 24506
rect 23175 24454 23187 24506
rect 23239 24454 23251 24506
rect 23303 24454 23315 24506
rect 23367 24454 34316 24506
rect 1104 24432 34316 24454
rect 1581 24395 1639 24401
rect 1581 24361 1593 24395
rect 1627 24392 1639 24395
rect 7558 24392 7564 24404
rect 1627 24364 7564 24392
rect 1627 24361 1639 24364
rect 1581 24355 1639 24361
rect 7558 24352 7564 24364
rect 7616 24352 7622 24404
rect 9030 24392 9036 24404
rect 7852 24364 9036 24392
rect 2777 24327 2835 24333
rect 2777 24293 2789 24327
rect 2823 24324 2835 24327
rect 2866 24324 2872 24336
rect 2823 24296 2872 24324
rect 2823 24293 2835 24296
rect 2777 24287 2835 24293
rect 2866 24284 2872 24296
rect 2924 24284 2930 24336
rect 6270 24324 6276 24336
rect 6183 24296 6276 24324
rect 6270 24284 6276 24296
rect 6328 24324 6334 24336
rect 7852 24324 7880 24364
rect 9030 24352 9036 24364
rect 9088 24392 9094 24404
rect 10594 24392 10600 24404
rect 9088 24364 10600 24392
rect 9088 24352 9094 24364
rect 10594 24352 10600 24364
rect 10652 24352 10658 24404
rect 10796 24364 11376 24392
rect 10796 24336 10824 24364
rect 6328 24296 7880 24324
rect 6328 24284 6334 24296
rect 7926 24284 7932 24336
rect 7984 24324 7990 24336
rect 8205 24327 8263 24333
rect 8205 24324 8217 24327
rect 7984 24296 8217 24324
rect 7984 24284 7990 24296
rect 8205 24293 8217 24296
rect 8251 24293 8263 24327
rect 8205 24287 8263 24293
rect 10778 24284 10784 24336
rect 10836 24284 10842 24336
rect 11238 24324 11244 24336
rect 11199 24296 11244 24324
rect 11238 24284 11244 24296
rect 11296 24284 11302 24336
rect 11348 24324 11376 24364
rect 11606 24352 11612 24404
rect 11664 24392 11670 24404
rect 11664 24364 12940 24392
rect 11664 24352 11670 24364
rect 11348 24296 12848 24324
rect 1394 24256 1400 24268
rect 1355 24228 1400 24256
rect 1394 24216 1400 24228
rect 1452 24216 1458 24268
rect 2130 24256 2136 24268
rect 2091 24228 2136 24256
rect 2130 24216 2136 24228
rect 2188 24216 2194 24268
rect 3145 24259 3203 24265
rect 3145 24225 3157 24259
rect 3191 24225 3203 24259
rect 3326 24256 3332 24268
rect 3287 24228 3332 24256
rect 3145 24219 3203 24225
rect 3160 24188 3188 24219
rect 3326 24216 3332 24228
rect 3384 24216 3390 24268
rect 4338 24216 4344 24268
rect 4396 24256 4402 24268
rect 4433 24259 4491 24265
rect 4433 24256 4445 24259
rect 4396 24228 4445 24256
rect 4396 24216 4402 24228
rect 4433 24225 4445 24228
rect 4479 24225 4491 24259
rect 5166 24256 5172 24268
rect 5127 24228 5172 24256
rect 4433 24219 4491 24225
rect 5166 24216 5172 24228
rect 5224 24216 5230 24268
rect 6181 24259 6239 24265
rect 6181 24225 6193 24259
rect 6227 24256 6239 24259
rect 6914 24256 6920 24268
rect 6227 24228 6920 24256
rect 6227 24225 6239 24228
rect 6181 24219 6239 24225
rect 6914 24216 6920 24228
rect 6972 24256 6978 24268
rect 6972 24228 7512 24256
rect 6972 24216 6978 24228
rect 4522 24188 4528 24200
rect 3160 24160 4528 24188
rect 4522 24148 4528 24160
rect 4580 24188 4586 24200
rect 5261 24191 5319 24197
rect 5261 24188 5273 24191
rect 4580 24160 5273 24188
rect 4580 24148 4586 24160
rect 5261 24157 5273 24160
rect 5307 24157 5319 24191
rect 5261 24151 5319 24157
rect 3145 24123 3203 24129
rect 3145 24089 3157 24123
rect 3191 24120 3203 24123
rect 3786 24120 3792 24132
rect 3191 24092 3792 24120
rect 3191 24089 3203 24092
rect 3145 24083 3203 24089
rect 3786 24080 3792 24092
rect 3844 24080 3850 24132
rect 4614 24120 4620 24132
rect 4575 24092 4620 24120
rect 4614 24080 4620 24092
rect 4672 24080 4678 24132
rect 1762 24012 1768 24064
rect 1820 24052 1826 24064
rect 2225 24055 2283 24061
rect 2225 24052 2237 24055
rect 1820 24024 2237 24052
rect 1820 24012 1826 24024
rect 2225 24021 2237 24024
rect 2271 24052 2283 24055
rect 2774 24052 2780 24064
rect 2271 24024 2780 24052
rect 2271 24021 2283 24024
rect 2225 24015 2283 24021
rect 2774 24012 2780 24024
rect 2832 24012 2838 24064
rect 7484 24052 7512 24228
rect 7558 24216 7564 24268
rect 7616 24256 7622 24268
rect 8021 24259 8079 24265
rect 8021 24256 8033 24259
rect 7616 24228 8033 24256
rect 7616 24216 7622 24228
rect 8021 24225 8033 24228
rect 8067 24225 8079 24259
rect 8021 24219 8079 24225
rect 8036 24188 8064 24219
rect 11790 24216 11796 24268
rect 11848 24256 11854 24268
rect 12161 24259 12219 24265
rect 12161 24256 12173 24259
rect 11848 24228 12173 24256
rect 11848 24216 11854 24228
rect 12161 24225 12173 24228
rect 12207 24225 12219 24259
rect 12161 24219 12219 24225
rect 11238 24188 11244 24200
rect 8036 24160 11244 24188
rect 11238 24148 11244 24160
rect 11296 24148 11302 24200
rect 11514 24188 11520 24200
rect 11475 24160 11520 24188
rect 11514 24148 11520 24160
rect 11572 24148 11578 24200
rect 12342 24148 12348 24200
rect 12400 24188 12406 24200
rect 12437 24191 12495 24197
rect 12437 24188 12449 24191
rect 12400 24160 12449 24188
rect 12400 24148 12406 24160
rect 12437 24157 12449 24160
rect 12483 24157 12495 24191
rect 12820 24188 12848 24296
rect 12912 24265 12940 24364
rect 12986 24352 12992 24404
rect 13044 24392 13050 24404
rect 18138 24392 18144 24404
rect 13044 24364 13089 24392
rect 18099 24364 18144 24392
rect 13044 24352 13050 24364
rect 18138 24352 18144 24364
rect 18196 24352 18202 24404
rect 18693 24395 18751 24401
rect 18693 24361 18705 24395
rect 18739 24361 18751 24395
rect 18693 24355 18751 24361
rect 20165 24395 20223 24401
rect 20165 24361 20177 24395
rect 20211 24392 20223 24395
rect 20438 24392 20444 24404
rect 20211 24364 20444 24392
rect 20211 24361 20223 24364
rect 20165 24355 20223 24361
rect 16298 24284 16304 24336
rect 16356 24324 16362 24336
rect 16356 24296 18184 24324
rect 16356 24284 16362 24296
rect 16408 24265 16436 24296
rect 12897 24259 12955 24265
rect 12897 24225 12909 24259
rect 12943 24225 12955 24259
rect 12897 24219 12955 24225
rect 16392 24259 16450 24265
rect 16392 24225 16404 24259
rect 16438 24225 16450 24259
rect 16392 24219 16450 24225
rect 16485 24259 16543 24265
rect 16485 24225 16497 24259
rect 16531 24225 16543 24259
rect 17126 24256 17132 24268
rect 17087 24228 17132 24256
rect 16485 24219 16543 24225
rect 14550 24188 14556 24200
rect 12820 24160 14556 24188
rect 12437 24151 12495 24157
rect 14550 24148 14556 24160
rect 14608 24148 14614 24200
rect 16500 24188 16528 24219
rect 17126 24216 17132 24228
rect 17184 24216 17190 24268
rect 18156 24265 18184 24296
rect 17957 24259 18015 24265
rect 17957 24256 17969 24259
rect 17512 24228 17969 24256
rect 17218 24188 17224 24200
rect 16500 24160 17224 24188
rect 17218 24148 17224 24160
rect 17276 24148 17282 24200
rect 8389 24123 8447 24129
rect 8389 24089 8401 24123
rect 8435 24120 8447 24123
rect 8662 24120 8668 24132
rect 8435 24092 8668 24120
rect 8435 24089 8447 24092
rect 8389 24083 8447 24089
rect 8662 24080 8668 24092
rect 8720 24080 8726 24132
rect 9950 24120 9956 24132
rect 8772 24092 9956 24120
rect 8772 24052 8800 24092
rect 9950 24080 9956 24092
rect 10008 24080 10014 24132
rect 11698 24080 11704 24132
rect 11756 24120 11762 24132
rect 15286 24120 15292 24132
rect 11756 24092 15292 24120
rect 11756 24080 11762 24092
rect 15286 24080 15292 24092
rect 15344 24080 15350 24132
rect 16114 24120 16120 24132
rect 16075 24092 16120 24120
rect 16114 24080 16120 24092
rect 16172 24080 16178 24132
rect 17512 24129 17540 24228
rect 17957 24225 17969 24228
rect 18003 24225 18015 24259
rect 17957 24219 18015 24225
rect 18141 24259 18199 24265
rect 18141 24225 18153 24259
rect 18187 24256 18199 24259
rect 18708 24256 18736 24355
rect 20438 24352 20444 24364
rect 20496 24352 20502 24404
rect 21082 24352 21088 24404
rect 21140 24392 21146 24404
rect 21140 24364 22416 24392
rect 21140 24352 21146 24364
rect 22388 24336 22416 24364
rect 22922 24352 22928 24404
rect 22980 24392 22986 24404
rect 23498 24395 23556 24401
rect 23498 24392 23510 24395
rect 22980 24364 23510 24392
rect 22980 24352 22986 24364
rect 23498 24361 23510 24364
rect 23544 24361 23556 24395
rect 23498 24355 23556 24361
rect 24305 24395 24363 24401
rect 24305 24361 24317 24395
rect 24351 24392 24363 24395
rect 25130 24392 25136 24404
rect 24351 24364 25136 24392
rect 24351 24361 24363 24364
rect 24305 24355 24363 24361
rect 25130 24352 25136 24364
rect 25188 24352 25194 24404
rect 27890 24392 27896 24404
rect 25240 24364 27896 24392
rect 18782 24284 18788 24336
rect 18840 24333 18846 24336
rect 18840 24327 18903 24333
rect 18840 24293 18857 24327
rect 18891 24293 18903 24327
rect 18840 24287 18903 24293
rect 19061 24327 19119 24333
rect 19061 24293 19073 24327
rect 19107 24293 19119 24327
rect 19061 24287 19119 24293
rect 18840 24284 18846 24287
rect 18187 24228 18736 24256
rect 19076 24256 19104 24287
rect 22370 24284 22376 24336
rect 22428 24284 22434 24336
rect 23014 24284 23020 24336
rect 23072 24324 23078 24336
rect 23293 24327 23351 24333
rect 23293 24324 23305 24327
rect 23072 24296 23305 24324
rect 23072 24284 23078 24296
rect 23293 24293 23305 24296
rect 23339 24324 23351 24327
rect 23339 24296 23796 24324
rect 23339 24293 23351 24296
rect 23293 24287 23351 24293
rect 19981 24259 20039 24265
rect 19981 24256 19993 24259
rect 19076 24228 19993 24256
rect 18187 24225 18199 24228
rect 18141 24219 18199 24225
rect 19981 24225 19993 24228
rect 20027 24256 20039 24259
rect 20027 24228 21496 24256
rect 20027 24225 20039 24228
rect 19981 24219 20039 24225
rect 20990 24188 20996 24200
rect 20951 24160 20996 24188
rect 20990 24148 20996 24160
rect 21048 24148 21054 24200
rect 21358 24188 21364 24200
rect 21319 24160 21364 24188
rect 21358 24148 21364 24160
rect 21416 24148 21422 24200
rect 21468 24188 21496 24228
rect 23768 24188 23796 24296
rect 23934 24284 23940 24336
rect 23992 24324 23998 24336
rect 23992 24296 24348 24324
rect 23992 24284 23998 24296
rect 23842 24216 23848 24268
rect 23900 24256 23906 24268
rect 24320 24265 24348 24296
rect 24121 24259 24179 24265
rect 24121 24256 24133 24259
rect 23900 24228 24133 24256
rect 23900 24216 23906 24228
rect 24121 24225 24133 24228
rect 24167 24225 24179 24259
rect 24121 24219 24179 24225
rect 24305 24259 24363 24265
rect 24305 24225 24317 24259
rect 24351 24225 24363 24259
rect 24305 24219 24363 24225
rect 25240 24188 25268 24364
rect 27890 24352 27896 24364
rect 27948 24352 27954 24404
rect 29178 24392 29184 24404
rect 29139 24364 29184 24392
rect 29178 24352 29184 24364
rect 29236 24352 29242 24404
rect 31202 24392 31208 24404
rect 31163 24364 31208 24392
rect 31202 24352 31208 24364
rect 31260 24352 31266 24404
rect 27154 24324 27160 24336
rect 27115 24296 27160 24324
rect 27154 24284 27160 24296
rect 27212 24284 27218 24336
rect 28442 24284 28448 24336
rect 28500 24324 28506 24336
rect 32122 24324 32128 24336
rect 28500 24296 29316 24324
rect 28500 24284 28506 24296
rect 25498 24256 25504 24268
rect 25459 24228 25504 24256
rect 25498 24216 25504 24228
rect 25556 24216 25562 24268
rect 25866 24256 25872 24268
rect 25827 24228 25872 24256
rect 25866 24216 25872 24228
rect 25924 24216 25930 24268
rect 25958 24216 25964 24268
rect 26016 24256 26022 24268
rect 29288 24265 29316 24296
rect 31864 24296 32128 24324
rect 29089 24259 29147 24265
rect 29089 24256 29101 24259
rect 26016 24228 26061 24256
rect 28290 24228 28488 24256
rect 26016 24216 26022 24228
rect 26878 24188 26884 24200
rect 21468 24160 23520 24188
rect 23768 24160 25268 24188
rect 26839 24160 26884 24188
rect 17497 24123 17555 24129
rect 17497 24089 17509 24123
rect 17543 24089 17555 24123
rect 17497 24083 17555 24089
rect 23492 24120 23520 24160
rect 26878 24148 26884 24160
rect 26936 24148 26942 24200
rect 28350 24188 28356 24200
rect 26988 24160 28356 24188
rect 26988 24120 27016 24160
rect 28350 24148 28356 24160
rect 28408 24148 28414 24200
rect 23492 24092 27016 24120
rect 28460 24120 28488 24228
rect 28644 24228 29101 24256
rect 28534 24148 28540 24200
rect 28592 24188 28598 24200
rect 28644 24197 28672 24228
rect 29089 24225 29101 24228
rect 29135 24225 29147 24259
rect 29089 24219 29147 24225
rect 29273 24259 29331 24265
rect 29273 24225 29285 24259
rect 29319 24225 29331 24259
rect 29273 24219 29331 24225
rect 30834 24216 30840 24268
rect 30892 24256 30898 24268
rect 31297 24259 31355 24265
rect 31297 24256 31309 24259
rect 30892 24228 31309 24256
rect 30892 24216 30898 24228
rect 31297 24225 31309 24228
rect 31343 24225 31355 24259
rect 31297 24219 31355 24225
rect 28629 24191 28687 24197
rect 28629 24188 28641 24191
rect 28592 24160 28641 24188
rect 28592 24148 28598 24160
rect 28629 24157 28641 24160
rect 28675 24157 28687 24191
rect 28629 24151 28687 24157
rect 31205 24191 31263 24197
rect 31205 24157 31217 24191
rect 31251 24188 31263 24191
rect 31386 24188 31392 24200
rect 31251 24160 31392 24188
rect 31251 24157 31263 24160
rect 31205 24151 31263 24157
rect 31386 24148 31392 24160
rect 31444 24148 31450 24200
rect 31754 24148 31760 24200
rect 31812 24188 31818 24200
rect 31864 24197 31892 24296
rect 32122 24284 32128 24296
rect 32180 24284 32186 24336
rect 32582 24284 32588 24336
rect 32640 24284 32646 24336
rect 31849 24191 31907 24197
rect 31849 24188 31861 24191
rect 31812 24160 31861 24188
rect 31812 24148 31818 24160
rect 31849 24157 31861 24160
rect 31895 24157 31907 24191
rect 31849 24151 31907 24157
rect 32125 24191 32183 24197
rect 32125 24157 32137 24191
rect 32171 24188 32183 24191
rect 32858 24188 32864 24200
rect 32171 24160 32864 24188
rect 32171 24157 32183 24160
rect 32125 24151 32183 24157
rect 32858 24148 32864 24160
rect 32916 24148 32922 24200
rect 29822 24120 29828 24132
rect 28460 24092 29828 24120
rect 7484 24024 8800 24052
rect 9769 24055 9827 24061
rect 9769 24021 9781 24055
rect 9815 24052 9827 24055
rect 11606 24052 11612 24064
rect 9815 24024 11612 24052
rect 9815 24021 9827 24024
rect 9769 24015 9827 24021
rect 11606 24012 11612 24024
rect 11664 24012 11670 24064
rect 12250 24052 12256 24064
rect 12211 24024 12256 24052
rect 12250 24012 12256 24024
rect 12308 24012 12314 24064
rect 12345 24055 12403 24061
rect 12345 24021 12357 24055
rect 12391 24052 12403 24055
rect 12894 24052 12900 24064
rect 12391 24024 12900 24052
rect 12391 24021 12403 24024
rect 12345 24015 12403 24021
rect 12894 24012 12900 24024
rect 12952 24012 12958 24064
rect 17954 24012 17960 24064
rect 18012 24052 18018 24064
rect 18877 24055 18935 24061
rect 18877 24052 18889 24055
rect 18012 24024 18889 24052
rect 18012 24012 18018 24024
rect 18877 24021 18889 24024
rect 18923 24021 18935 24055
rect 18877 24015 18935 24021
rect 22787 24055 22845 24061
rect 22787 24021 22799 24055
rect 22833 24052 22845 24055
rect 23014 24052 23020 24064
rect 22833 24024 23020 24052
rect 22833 24021 22845 24024
rect 22787 24015 22845 24021
rect 23014 24012 23020 24024
rect 23072 24012 23078 24064
rect 23492 24061 23520 24092
rect 29822 24080 29828 24092
rect 29880 24080 29886 24132
rect 23477 24055 23535 24061
rect 23477 24021 23489 24055
rect 23523 24021 23535 24055
rect 23658 24052 23664 24064
rect 23619 24024 23664 24052
rect 23477 24015 23535 24021
rect 23658 24012 23664 24024
rect 23716 24012 23722 24064
rect 24394 24012 24400 24064
rect 24452 24052 24458 24064
rect 25317 24055 25375 24061
rect 25317 24052 25329 24055
rect 24452 24024 25329 24052
rect 24452 24012 24458 24024
rect 25317 24021 25329 24024
rect 25363 24021 25375 24055
rect 30742 24052 30748 24064
rect 30703 24024 30748 24052
rect 25317 24015 25375 24021
rect 30742 24012 30748 24024
rect 30800 24012 30806 24064
rect 33594 24052 33600 24064
rect 33555 24024 33600 24052
rect 33594 24012 33600 24024
rect 33652 24012 33658 24064
rect 1104 23962 34316 23984
rect 1104 23910 6517 23962
rect 6569 23910 6581 23962
rect 6633 23910 6645 23962
rect 6697 23910 6709 23962
rect 6761 23910 17588 23962
rect 17640 23910 17652 23962
rect 17704 23910 17716 23962
rect 17768 23910 17780 23962
rect 17832 23910 28658 23962
rect 28710 23910 28722 23962
rect 28774 23910 28786 23962
rect 28838 23910 28850 23962
rect 28902 23910 34316 23962
rect 1104 23888 34316 23910
rect 2685 23851 2743 23857
rect 2685 23817 2697 23851
rect 2731 23848 2743 23851
rect 2958 23848 2964 23860
rect 2731 23820 2964 23848
rect 2731 23817 2743 23820
rect 2685 23811 2743 23817
rect 2958 23808 2964 23820
rect 3016 23808 3022 23860
rect 8846 23808 8852 23860
rect 8904 23848 8910 23860
rect 9217 23851 9275 23857
rect 9217 23848 9229 23851
rect 8904 23820 9229 23848
rect 8904 23808 8910 23820
rect 9217 23817 9229 23820
rect 9263 23817 9275 23851
rect 9217 23811 9275 23817
rect 9582 23808 9588 23860
rect 9640 23848 9646 23860
rect 10505 23851 10563 23857
rect 10505 23848 10517 23851
rect 9640 23820 10517 23848
rect 9640 23808 9646 23820
rect 10505 23817 10517 23820
rect 10551 23817 10563 23851
rect 10505 23811 10563 23817
rect 10594 23808 10600 23860
rect 10652 23848 10658 23860
rect 11698 23848 11704 23860
rect 10652 23820 11704 23848
rect 10652 23808 10658 23820
rect 11698 23808 11704 23820
rect 11756 23808 11762 23860
rect 12342 23848 12348 23860
rect 12303 23820 12348 23848
rect 12342 23808 12348 23820
rect 12400 23808 12406 23860
rect 19426 23848 19432 23860
rect 19387 23820 19432 23848
rect 19426 23808 19432 23820
rect 19484 23808 19490 23860
rect 25317 23851 25375 23857
rect 25317 23817 25329 23851
rect 25363 23848 25375 23851
rect 26878 23848 26884 23860
rect 25363 23820 26884 23848
rect 25363 23817 25375 23820
rect 25317 23811 25375 23817
rect 26878 23808 26884 23820
rect 26936 23808 26942 23860
rect 3513 23783 3571 23789
rect 3513 23749 3525 23783
rect 3559 23780 3571 23783
rect 4338 23780 4344 23792
rect 3559 23752 4344 23780
rect 3559 23749 3571 23752
rect 3513 23743 3571 23749
rect 4338 23740 4344 23752
rect 4396 23740 4402 23792
rect 9861 23783 9919 23789
rect 9861 23780 9873 23783
rect 8036 23752 9873 23780
rect 4430 23712 4436 23724
rect 4391 23684 4436 23712
rect 4430 23672 4436 23684
rect 4488 23672 4494 23724
rect 4614 23672 4620 23724
rect 4672 23712 4678 23724
rect 8036 23721 8064 23752
rect 9861 23749 9873 23752
rect 9907 23749 9919 23783
rect 9861 23743 9919 23749
rect 11514 23740 11520 23792
rect 11572 23780 11578 23792
rect 29454 23780 29460 23792
rect 11572 23752 12756 23780
rect 29415 23752 29460 23780
rect 11572 23740 11578 23752
rect 4985 23715 5043 23721
rect 4985 23712 4997 23715
rect 4672 23684 4997 23712
rect 4672 23672 4678 23684
rect 4985 23681 4997 23684
rect 5031 23681 5043 23715
rect 4985 23675 5043 23681
rect 8021 23715 8079 23721
rect 8021 23681 8033 23715
rect 8067 23681 8079 23715
rect 8021 23675 8079 23681
rect 8205 23715 8263 23721
rect 8205 23681 8217 23715
rect 8251 23712 8263 23715
rect 8757 23715 8815 23721
rect 8757 23712 8769 23715
rect 8251 23684 8769 23712
rect 8251 23681 8263 23684
rect 8205 23675 8263 23681
rect 8757 23681 8769 23684
rect 8803 23681 8815 23715
rect 9122 23712 9128 23724
rect 8757 23675 8815 23681
rect 8956 23684 9128 23712
rect 2777 23647 2835 23653
rect 2777 23613 2789 23647
rect 2823 23613 2835 23647
rect 2777 23607 2835 23613
rect 4801 23647 4859 23653
rect 4801 23613 4813 23647
rect 4847 23644 4859 23647
rect 4890 23644 4896 23656
rect 4847 23616 4896 23644
rect 4847 23613 4859 23616
rect 4801 23607 4859 23613
rect 2792 23576 2820 23607
rect 4890 23604 4896 23616
rect 4948 23604 4954 23656
rect 5258 23604 5264 23656
rect 5316 23644 5322 23656
rect 5353 23647 5411 23653
rect 5353 23644 5365 23647
rect 5316 23616 5365 23644
rect 5316 23604 5322 23616
rect 5353 23613 5365 23616
rect 5399 23613 5411 23647
rect 5353 23607 5411 23613
rect 5813 23647 5871 23653
rect 5813 23613 5825 23647
rect 5859 23644 5871 23647
rect 6914 23644 6920 23656
rect 5859 23616 6920 23644
rect 5859 23613 5871 23616
rect 5813 23607 5871 23613
rect 6914 23604 6920 23616
rect 6972 23604 6978 23656
rect 8956 23653 8984 23684
rect 9122 23672 9128 23684
rect 9180 23672 9186 23724
rect 10226 23712 10232 23724
rect 9324 23684 10232 23712
rect 8297 23647 8355 23653
rect 8297 23613 8309 23647
rect 8343 23613 8355 23647
rect 8297 23607 8355 23613
rect 8941 23647 8999 23653
rect 8941 23613 8953 23647
rect 8987 23613 8999 23647
rect 8941 23607 8999 23613
rect 9033 23647 9091 23653
rect 9033 23613 9045 23647
rect 9079 23644 9091 23647
rect 9214 23644 9220 23656
rect 9079 23616 9220 23644
rect 9079 23613 9091 23616
rect 9033 23607 9091 23613
rect 3326 23576 3332 23588
rect 2792 23548 3332 23576
rect 3326 23536 3332 23548
rect 3384 23536 3390 23588
rect 8312 23576 8340 23607
rect 9214 23604 9220 23616
rect 9272 23604 9278 23656
rect 9324 23653 9352 23684
rect 10226 23672 10232 23684
rect 10284 23672 10290 23724
rect 10318 23672 10324 23724
rect 10376 23712 10382 23724
rect 12434 23712 12440 23724
rect 10376 23684 10640 23712
rect 10376 23672 10382 23684
rect 9309 23647 9367 23653
rect 9309 23613 9321 23647
rect 9355 23613 9367 23647
rect 9766 23644 9772 23656
rect 9727 23616 9772 23644
rect 9309 23607 9367 23613
rect 9766 23604 9772 23616
rect 9824 23604 9830 23656
rect 9950 23644 9956 23656
rect 9911 23616 9956 23644
rect 9950 23604 9956 23616
rect 10008 23604 10014 23656
rect 10612 23653 10640 23684
rect 12268 23684 12440 23712
rect 10413 23647 10471 23653
rect 10413 23613 10425 23647
rect 10459 23613 10471 23647
rect 10413 23607 10471 23613
rect 10597 23647 10655 23653
rect 10597 23613 10609 23647
rect 10643 23613 10655 23647
rect 10597 23607 10655 23613
rect 9784 23576 9812 23604
rect 8312 23548 9812 23576
rect 8021 23511 8079 23517
rect 8021 23477 8033 23511
rect 8067 23508 8079 23511
rect 8386 23508 8392 23520
rect 8067 23480 8392 23508
rect 8067 23477 8079 23480
rect 8021 23471 8079 23477
rect 8386 23468 8392 23480
rect 8444 23468 8450 23520
rect 8478 23468 8484 23520
rect 8536 23508 8542 23520
rect 10428 23508 10456 23607
rect 11422 23604 11428 23656
rect 11480 23644 11486 23656
rect 12268 23653 12296 23684
rect 12434 23672 12440 23684
rect 12492 23672 12498 23724
rect 12161 23647 12219 23653
rect 12161 23644 12173 23647
rect 11480 23616 12173 23644
rect 11480 23604 11486 23616
rect 12161 23613 12173 23616
rect 12207 23613 12219 23647
rect 12161 23607 12219 23613
rect 12253 23647 12311 23653
rect 12253 23613 12265 23647
rect 12299 23613 12311 23647
rect 12728 23644 12756 23752
rect 29454 23740 29460 23752
rect 29512 23740 29518 23792
rect 12894 23672 12900 23724
rect 12952 23712 12958 23724
rect 13449 23715 13507 23721
rect 13449 23712 13461 23715
rect 12952 23684 13461 23712
rect 12952 23672 12958 23684
rect 13449 23681 13461 23684
rect 13495 23681 13507 23715
rect 25222 23712 25228 23724
rect 13449 23675 13507 23681
rect 22940 23684 25228 23712
rect 13173 23647 13231 23653
rect 13173 23644 13185 23647
rect 12728 23616 13185 23644
rect 12253 23607 12311 23613
rect 13173 23613 13185 23616
rect 13219 23613 13231 23647
rect 13173 23607 13231 23613
rect 12437 23579 12495 23585
rect 12437 23545 12449 23579
rect 12483 23576 12495 23579
rect 12618 23576 12624 23588
rect 12483 23548 12624 23576
rect 12483 23545 12495 23548
rect 12437 23539 12495 23545
rect 12618 23536 12624 23548
rect 12676 23536 12682 23588
rect 13188 23576 13216 23607
rect 14550 23604 14556 23656
rect 14608 23644 14614 23656
rect 15470 23644 15476 23656
rect 14608 23616 15476 23644
rect 14608 23604 14614 23616
rect 15470 23604 15476 23616
rect 15528 23604 15534 23656
rect 22940 23653 22968 23684
rect 19705 23647 19763 23653
rect 19705 23613 19717 23647
rect 19751 23644 19763 23647
rect 22925 23647 22983 23653
rect 19751 23616 22094 23644
rect 19751 23613 19763 23616
rect 19705 23607 19763 23613
rect 13722 23576 13728 23588
rect 13188 23548 13728 23576
rect 13722 23536 13728 23548
rect 13780 23536 13786 23588
rect 19429 23579 19487 23585
rect 19429 23545 19441 23579
rect 19475 23576 19487 23579
rect 20622 23576 20628 23588
rect 19475 23548 20628 23576
rect 19475 23545 19487 23548
rect 19429 23539 19487 23545
rect 20622 23536 20628 23548
rect 20680 23536 20686 23588
rect 22066 23576 22094 23616
rect 22925 23613 22937 23647
rect 22971 23613 22983 23647
rect 22925 23607 22983 23613
rect 23385 23647 23443 23653
rect 23385 23613 23397 23647
rect 23431 23644 23443 23647
rect 23474 23644 23480 23656
rect 23431 23616 23480 23644
rect 23431 23613 23443 23616
rect 23385 23607 23443 23613
rect 23474 23604 23480 23616
rect 23532 23604 23538 23656
rect 23842 23644 23848 23656
rect 23803 23616 23848 23644
rect 23842 23604 23848 23616
rect 23900 23604 23906 23656
rect 24213 23647 24271 23653
rect 24213 23613 24225 23647
rect 24259 23644 24271 23647
rect 24394 23644 24400 23656
rect 24259 23616 24400 23644
rect 24259 23613 24271 23616
rect 24213 23607 24271 23613
rect 24394 23604 24400 23616
rect 24452 23604 24458 23656
rect 25148 23653 25176 23684
rect 25222 23672 25228 23684
rect 25280 23672 25286 23724
rect 28442 23712 28448 23724
rect 28368 23684 28448 23712
rect 28368 23653 28396 23684
rect 28442 23672 28448 23684
rect 28500 23672 28506 23724
rect 30742 23712 30748 23724
rect 30130 23684 30748 23712
rect 30742 23672 30748 23684
rect 30800 23672 30806 23724
rect 30837 23715 30895 23721
rect 30837 23681 30849 23715
rect 30883 23712 30895 23715
rect 30883 23684 31892 23712
rect 30883 23681 30895 23684
rect 30837 23675 30895 23681
rect 25133 23647 25191 23653
rect 25133 23613 25145 23647
rect 25179 23613 25191 23647
rect 25133 23607 25191 23613
rect 25409 23647 25467 23653
rect 25409 23613 25421 23647
rect 25455 23613 25467 23647
rect 25409 23607 25467 23613
rect 28353 23647 28411 23653
rect 28353 23613 28365 23647
rect 28399 23613 28411 23647
rect 28534 23644 28540 23656
rect 28495 23616 28540 23644
rect 28353 23607 28411 23613
rect 23566 23576 23572 23588
rect 22066 23548 23572 23576
rect 23566 23536 23572 23548
rect 23624 23536 23630 23588
rect 24302 23576 24308 23588
rect 24263 23548 24308 23576
rect 24302 23536 24308 23548
rect 24360 23536 24366 23588
rect 24486 23536 24492 23588
rect 24544 23576 24550 23588
rect 25424 23576 25452 23607
rect 28534 23604 28540 23616
rect 28592 23604 28598 23656
rect 29638 23644 29644 23656
rect 29599 23616 29644 23644
rect 29638 23604 29644 23616
rect 29696 23604 29702 23656
rect 30466 23644 30472 23656
rect 30427 23616 30472 23644
rect 30466 23604 30472 23616
rect 30524 23604 30530 23656
rect 30760 23644 30788 23672
rect 31864 23656 31892 23684
rect 31573 23647 31631 23653
rect 31573 23644 31585 23647
rect 30760 23616 31585 23644
rect 31573 23613 31585 23616
rect 31619 23613 31631 23647
rect 31846 23644 31852 23656
rect 31807 23616 31852 23644
rect 31573 23607 31631 23613
rect 31846 23604 31852 23616
rect 31904 23604 31910 23656
rect 24544 23548 25452 23576
rect 24544 23536 24550 23548
rect 25498 23536 25504 23588
rect 25556 23576 25562 23588
rect 25654 23579 25712 23585
rect 25654 23576 25666 23579
rect 25556 23548 25666 23576
rect 25556 23536 25562 23548
rect 25654 23545 25666 23548
rect 25700 23545 25712 23579
rect 25654 23539 25712 23545
rect 8536 23480 10456 23508
rect 8536 23468 8542 23480
rect 13262 23468 13268 23520
rect 13320 23508 13326 23520
rect 13630 23508 13636 23520
rect 13320 23480 13636 23508
rect 13320 23468 13326 23480
rect 13630 23468 13636 23480
rect 13688 23508 13694 23520
rect 14921 23511 14979 23517
rect 14921 23508 14933 23511
rect 13688 23480 14933 23508
rect 13688 23468 13694 23480
rect 14921 23477 14933 23480
rect 14967 23477 14979 23511
rect 19610 23508 19616 23520
rect 19571 23480 19616 23508
rect 14921 23471 14979 23477
rect 19610 23468 19616 23480
rect 19668 23468 19674 23520
rect 20162 23468 20168 23520
rect 20220 23508 20226 23520
rect 20990 23508 20996 23520
rect 20220 23480 20996 23508
rect 20220 23468 20226 23480
rect 20990 23468 20996 23480
rect 21048 23508 21054 23520
rect 22741 23511 22799 23517
rect 22741 23508 22753 23511
rect 21048 23480 22753 23508
rect 21048 23468 21054 23480
rect 22741 23477 22753 23480
rect 22787 23508 22799 23511
rect 24504 23508 24532 23536
rect 26786 23508 26792 23520
rect 22787 23480 24532 23508
rect 26747 23480 26792 23508
rect 22787 23477 22799 23480
rect 22741 23471 22799 23477
rect 26786 23468 26792 23480
rect 26844 23468 26850 23520
rect 28166 23508 28172 23520
rect 28127 23480 28172 23508
rect 28166 23468 28172 23480
rect 28224 23468 28230 23520
rect 30484 23508 30512 23604
rect 30650 23536 30656 23588
rect 30708 23576 30714 23588
rect 31389 23579 31447 23585
rect 31389 23576 31401 23579
rect 30708 23548 31401 23576
rect 30708 23536 30714 23548
rect 31389 23545 31401 23548
rect 31435 23545 31447 23579
rect 31389 23539 31447 23545
rect 31757 23511 31815 23517
rect 31757 23508 31769 23511
rect 30484 23480 31769 23508
rect 31757 23477 31769 23480
rect 31803 23477 31815 23511
rect 31757 23471 31815 23477
rect 1104 23418 34316 23440
rect 1104 23366 12052 23418
rect 12104 23366 12116 23418
rect 12168 23366 12180 23418
rect 12232 23366 12244 23418
rect 12296 23366 23123 23418
rect 23175 23366 23187 23418
rect 23239 23366 23251 23418
rect 23303 23366 23315 23418
rect 23367 23366 34316 23418
rect 1104 23344 34316 23366
rect 9122 23264 9128 23316
rect 9180 23304 9186 23316
rect 9950 23304 9956 23316
rect 9180 23276 9956 23304
rect 9180 23264 9186 23276
rect 9950 23264 9956 23276
rect 10008 23304 10014 23316
rect 11054 23304 11060 23316
rect 10008 23276 11060 23304
rect 10008 23264 10014 23276
rect 2682 23196 2688 23248
rect 2740 23196 2746 23248
rect 5166 23196 5172 23248
rect 5224 23236 5230 23248
rect 5224 23208 7696 23236
rect 5224 23196 5230 23208
rect 2958 23128 2964 23180
rect 3016 23168 3022 23180
rect 5920 23177 5948 23208
rect 5077 23171 5135 23177
rect 5077 23168 5089 23171
rect 3016 23140 5089 23168
rect 3016 23128 3022 23140
rect 5077 23137 5089 23140
rect 5123 23137 5135 23171
rect 5077 23131 5135 23137
rect 5905 23171 5963 23177
rect 5905 23137 5917 23171
rect 5951 23137 5963 23171
rect 7098 23168 7104 23180
rect 7059 23140 7104 23168
rect 5905 23131 5963 23137
rect 7098 23128 7104 23140
rect 7156 23128 7162 23180
rect 7668 23177 7696 23208
rect 9766 23196 9772 23248
rect 9824 23236 9830 23248
rect 10137 23239 10195 23245
rect 10137 23236 10149 23239
rect 9824 23208 10149 23236
rect 9824 23196 9830 23208
rect 10137 23205 10149 23208
rect 10183 23205 10195 23239
rect 10137 23199 10195 23205
rect 7653 23171 7711 23177
rect 7653 23137 7665 23171
rect 7699 23137 7711 23171
rect 10042 23168 10048 23180
rect 10003 23140 10048 23168
rect 7653 23131 7711 23137
rect 10042 23128 10048 23140
rect 10100 23128 10106 23180
rect 10796 23177 10824 23276
rect 11054 23264 11060 23276
rect 11112 23264 11118 23316
rect 11882 23264 11888 23316
rect 11940 23304 11946 23316
rect 11977 23307 12035 23313
rect 11977 23304 11989 23307
rect 11940 23276 11989 23304
rect 11940 23264 11946 23276
rect 11977 23273 11989 23276
rect 12023 23273 12035 23307
rect 11977 23267 12035 23273
rect 14182 23264 14188 23316
rect 14240 23304 14246 23316
rect 14734 23304 14740 23316
rect 14240 23276 14740 23304
rect 14240 23264 14246 23276
rect 14734 23264 14740 23276
rect 14792 23304 14798 23316
rect 14829 23307 14887 23313
rect 14829 23304 14841 23307
rect 14792 23276 14841 23304
rect 14792 23264 14798 23276
rect 14829 23273 14841 23276
rect 14875 23273 14887 23307
rect 14829 23267 14887 23273
rect 17221 23307 17279 23313
rect 17221 23273 17233 23307
rect 17267 23304 17279 23307
rect 17402 23304 17408 23316
rect 17267 23276 17408 23304
rect 17267 23273 17279 23276
rect 17221 23267 17279 23273
rect 17402 23264 17408 23276
rect 17460 23264 17466 23316
rect 17865 23307 17923 23313
rect 17865 23273 17877 23307
rect 17911 23304 17923 23307
rect 17954 23304 17960 23316
rect 17911 23276 17960 23304
rect 17911 23273 17923 23276
rect 17865 23267 17923 23273
rect 11422 23196 11428 23248
rect 11480 23236 11486 23248
rect 12069 23239 12127 23245
rect 11480 23208 12020 23236
rect 11480 23196 11486 23208
rect 10321 23171 10379 23177
rect 10321 23137 10333 23171
rect 10367 23137 10379 23171
rect 10321 23131 10379 23137
rect 10597 23171 10655 23177
rect 10597 23137 10609 23171
rect 10643 23137 10655 23171
rect 10597 23131 10655 23137
rect 10781 23171 10839 23177
rect 10781 23137 10793 23171
rect 10827 23137 10839 23171
rect 10781 23131 10839 23137
rect 1394 23100 1400 23112
rect 1355 23072 1400 23100
rect 1394 23060 1400 23072
rect 1452 23060 1458 23112
rect 1673 23103 1731 23109
rect 1673 23069 1685 23103
rect 1719 23100 1731 23103
rect 4154 23100 4160 23112
rect 1719 23072 4160 23100
rect 1719 23069 1731 23072
rect 1673 23063 1731 23069
rect 4154 23060 4160 23072
rect 4212 23060 4218 23112
rect 5350 23100 5356 23112
rect 5311 23072 5356 23100
rect 5350 23060 5356 23072
rect 5408 23060 5414 23112
rect 5629 23103 5687 23109
rect 5629 23069 5641 23103
rect 5675 23100 5687 23103
rect 5810 23100 5816 23112
rect 5675 23072 5816 23100
rect 5675 23069 5687 23072
rect 5629 23063 5687 23069
rect 5810 23060 5816 23072
rect 5868 23060 5874 23112
rect 9306 23060 9312 23112
rect 9364 23100 9370 23112
rect 10336 23100 10364 23131
rect 9364 23072 10364 23100
rect 10612 23100 10640 23131
rect 11238 23128 11244 23180
rect 11296 23168 11302 23180
rect 11885 23171 11943 23177
rect 11885 23168 11897 23171
rect 11296 23140 11897 23168
rect 11296 23128 11302 23140
rect 11885 23137 11897 23140
rect 11931 23137 11943 23171
rect 11992 23168 12020 23208
rect 12069 23205 12081 23239
rect 12115 23236 12127 23239
rect 12434 23236 12440 23248
rect 12115 23208 12440 23236
rect 12115 23205 12127 23208
rect 12069 23199 12127 23205
rect 12434 23196 12440 23208
rect 12492 23196 12498 23248
rect 16114 23245 16120 23248
rect 16108 23236 16120 23245
rect 16075 23208 16120 23236
rect 16108 23199 16120 23208
rect 16114 23196 16120 23199
rect 16172 23196 16178 23248
rect 16298 23196 16304 23248
rect 16356 23196 16362 23248
rect 16666 23196 16672 23248
rect 16724 23236 16730 23248
rect 17880 23236 17908 23267
rect 17954 23264 17960 23276
rect 18012 23264 18018 23316
rect 20901 23307 20959 23313
rect 20901 23273 20913 23307
rect 20947 23304 20959 23307
rect 21358 23304 21364 23316
rect 20947 23276 21364 23304
rect 20947 23273 20959 23276
rect 20901 23267 20959 23273
rect 21358 23264 21364 23276
rect 21416 23264 21422 23316
rect 25317 23307 25375 23313
rect 25317 23273 25329 23307
rect 25363 23304 25375 23307
rect 25498 23304 25504 23316
rect 25363 23276 25504 23304
rect 25363 23273 25375 23276
rect 25317 23267 25375 23273
rect 25498 23264 25504 23276
rect 25556 23264 25562 23316
rect 28442 23304 28448 23316
rect 25700 23276 28448 23304
rect 16724 23208 17908 23236
rect 18969 23239 19027 23245
rect 16724 23196 16730 23208
rect 18969 23205 18981 23239
rect 19015 23236 19027 23239
rect 19610 23236 19616 23248
rect 19015 23208 19616 23236
rect 19015 23205 19027 23208
rect 18969 23199 19027 23205
rect 19610 23196 19616 23208
rect 19668 23196 19674 23248
rect 20533 23239 20591 23245
rect 20533 23205 20545 23239
rect 20579 23236 20591 23239
rect 23014 23236 23020 23248
rect 20579 23208 23020 23236
rect 20579 23205 20591 23208
rect 20533 23199 20591 23205
rect 23014 23196 23020 23208
rect 23072 23196 23078 23248
rect 23474 23196 23480 23248
rect 23532 23245 23538 23248
rect 23532 23239 23595 23245
rect 23532 23205 23549 23239
rect 23583 23205 23595 23239
rect 23532 23199 23595 23205
rect 23753 23239 23811 23245
rect 23753 23205 23765 23239
rect 23799 23236 23811 23239
rect 24394 23236 24400 23248
rect 23799 23208 24400 23236
rect 23799 23205 23811 23208
rect 23753 23199 23811 23205
rect 23532 23196 23538 23199
rect 24394 23196 24400 23208
rect 24452 23196 24458 23248
rect 25130 23196 25136 23248
rect 25188 23236 25194 23248
rect 25700 23236 25728 23276
rect 28442 23264 28448 23276
rect 28500 23304 28506 23316
rect 28721 23307 28779 23313
rect 28721 23304 28733 23307
rect 28500 23276 28733 23304
rect 28500 23264 28506 23276
rect 28721 23273 28733 23276
rect 28767 23273 28779 23307
rect 31754 23304 31760 23316
rect 28721 23267 28779 23273
rect 30668 23276 31760 23304
rect 25188 23208 25728 23236
rect 25777 23239 25835 23245
rect 25188 23196 25194 23208
rect 25777 23205 25789 23239
rect 25823 23236 25835 23239
rect 26786 23236 26792 23248
rect 25823 23208 26792 23236
rect 25823 23205 25835 23208
rect 25777 23199 25835 23205
rect 26786 23196 26792 23208
rect 26844 23196 26850 23248
rect 28258 23196 28264 23248
rect 28316 23236 28322 23248
rect 28316 23208 28856 23236
rect 28316 23196 28322 23208
rect 12161 23171 12219 23177
rect 12161 23168 12173 23171
rect 11992 23140 12173 23168
rect 11885 23131 11943 23137
rect 12161 23137 12173 23140
rect 12207 23137 12219 23171
rect 12161 23131 12219 23137
rect 12621 23171 12679 23177
rect 12621 23137 12633 23171
rect 12667 23137 12679 23171
rect 12621 23131 12679 23137
rect 12636 23100 12664 23131
rect 12710 23128 12716 23180
rect 12768 23168 12774 23180
rect 12805 23171 12863 23177
rect 12805 23168 12817 23171
rect 12768 23140 12817 23168
rect 12768 23128 12774 23140
rect 12805 23137 12817 23140
rect 12851 23137 12863 23171
rect 12805 23131 12863 23137
rect 14921 23171 14979 23177
rect 14921 23137 14933 23171
rect 14967 23168 14979 23171
rect 15010 23168 15016 23180
rect 14967 23140 15016 23168
rect 14967 23137 14979 23140
rect 14921 23131 14979 23137
rect 15010 23128 15016 23140
rect 15068 23128 15074 23180
rect 15841 23171 15899 23177
rect 15841 23137 15853 23171
rect 15887 23168 15899 23171
rect 16316 23168 16344 23196
rect 15887 23140 16344 23168
rect 15887 23137 15899 23140
rect 15841 23131 15899 23137
rect 17218 23128 17224 23180
rect 17276 23168 17282 23180
rect 17681 23171 17739 23177
rect 17681 23168 17693 23171
rect 17276 23140 17693 23168
rect 17276 23128 17282 23140
rect 17681 23137 17693 23140
rect 17727 23168 17739 23171
rect 18690 23168 18696 23180
rect 17727 23140 18696 23168
rect 17727 23137 17739 23140
rect 17681 23131 17739 23137
rect 18690 23128 18696 23140
rect 18748 23128 18754 23180
rect 18785 23171 18843 23177
rect 18785 23137 18797 23171
rect 18831 23137 18843 23171
rect 18785 23131 18843 23137
rect 19061 23171 19119 23177
rect 19061 23137 19073 23171
rect 19107 23168 19119 23171
rect 19334 23168 19340 23180
rect 19107 23140 19340 23168
rect 19107 23137 19119 23140
rect 19061 23131 19119 23137
rect 14366 23100 14372 23112
rect 10612 23072 14372 23100
rect 9364 23060 9370 23072
rect 10888 23044 10916 23072
rect 14366 23060 14372 23072
rect 14424 23060 14430 23112
rect 18800 23100 18828 23131
rect 19334 23128 19340 23140
rect 19392 23128 19398 23180
rect 20349 23171 20407 23177
rect 20349 23137 20361 23171
rect 20395 23137 20407 23171
rect 20349 23131 20407 23137
rect 19518 23100 19524 23112
rect 18800 23072 19524 23100
rect 19518 23060 19524 23072
rect 19576 23060 19582 23112
rect 20364 23100 20392 23131
rect 20438 23128 20444 23180
rect 20496 23168 20502 23180
rect 20625 23171 20683 23177
rect 20625 23168 20637 23171
rect 20496 23140 20637 23168
rect 20496 23128 20502 23140
rect 20625 23137 20637 23140
rect 20671 23137 20683 23171
rect 20625 23131 20683 23137
rect 20714 23128 20720 23180
rect 20772 23168 20778 23180
rect 22370 23168 22376 23180
rect 20772 23140 20817 23168
rect 22283 23140 22376 23168
rect 20772 23128 20778 23140
rect 22370 23128 22376 23140
rect 22428 23168 22434 23180
rect 24762 23168 24768 23180
rect 22428 23140 24768 23168
rect 22428 23128 22434 23140
rect 24762 23128 24768 23140
rect 24820 23128 24826 23180
rect 25685 23171 25743 23177
rect 25685 23137 25697 23171
rect 25731 23168 25743 23171
rect 25958 23168 25964 23180
rect 25731 23140 25964 23168
rect 25731 23137 25743 23140
rect 25685 23131 25743 23137
rect 25958 23128 25964 23140
rect 26016 23128 26022 23180
rect 27801 23171 27859 23177
rect 27801 23137 27813 23171
rect 27847 23168 27859 23171
rect 28166 23168 28172 23180
rect 27847 23140 28172 23168
rect 27847 23137 27859 23140
rect 27801 23131 27859 23137
rect 28166 23128 28172 23140
rect 28224 23128 28230 23180
rect 28828 23168 28856 23208
rect 28828 23140 28948 23168
rect 20806 23100 20812 23112
rect 20364 23072 20812 23100
rect 20806 23060 20812 23072
rect 20864 23060 20870 23112
rect 21726 23100 21732 23112
rect 21687 23072 21732 23100
rect 21726 23060 21732 23072
rect 21784 23060 21790 23112
rect 25774 23060 25780 23112
rect 25832 23100 25838 23112
rect 28920 23109 28948 23140
rect 29362 23128 29368 23180
rect 29420 23168 29426 23180
rect 30668 23177 30696 23276
rect 31754 23264 31760 23276
rect 31812 23264 31818 23316
rect 32858 23304 32864 23316
rect 32819 23276 32864 23304
rect 32858 23264 32864 23276
rect 32916 23264 32922 23316
rect 32950 23264 32956 23316
rect 33008 23304 33014 23316
rect 33229 23307 33287 23313
rect 33229 23304 33241 23307
rect 33008 23276 33241 23304
rect 33008 23264 33014 23276
rect 33229 23273 33241 23276
rect 33275 23304 33287 23307
rect 33594 23304 33600 23316
rect 33275 23276 33600 23304
rect 33275 23273 33287 23276
rect 33229 23267 33287 23273
rect 33594 23264 33600 23276
rect 33652 23264 33658 23316
rect 30653 23171 30711 23177
rect 30653 23168 30665 23171
rect 29420 23140 30665 23168
rect 29420 23128 29426 23140
rect 30653 23137 30665 23140
rect 30699 23137 30711 23171
rect 32582 23168 32588 23180
rect 32062 23140 32588 23168
rect 30653 23131 30711 23137
rect 32582 23128 32588 23140
rect 32640 23128 32646 23180
rect 25869 23103 25927 23109
rect 25869 23100 25881 23103
rect 25832 23072 25881 23100
rect 25832 23060 25838 23072
rect 25869 23069 25881 23072
rect 25915 23069 25927 23103
rect 25869 23063 25927 23069
rect 28813 23103 28871 23109
rect 28813 23069 28825 23103
rect 28859 23069 28871 23103
rect 28813 23063 28871 23069
rect 28905 23103 28963 23109
rect 28905 23069 28917 23103
rect 28951 23069 28963 23103
rect 30926 23100 30932 23112
rect 30887 23072 30932 23100
rect 28905 23063 28963 23069
rect 4801 23035 4859 23041
rect 4801 23001 4813 23035
rect 4847 23032 4859 23035
rect 4890 23032 4896 23044
rect 4847 23004 4896 23032
rect 4847 23001 4859 23004
rect 4801 22995 4859 23001
rect 4890 22992 4896 23004
rect 4948 22992 4954 23044
rect 8018 23032 8024 23044
rect 7979 23004 8024 23032
rect 8018 22992 8024 23004
rect 8076 23032 8082 23044
rect 8294 23032 8300 23044
rect 8076 23004 8300 23032
rect 8076 22992 8082 23004
rect 8294 22992 8300 23004
rect 8352 22992 8358 23044
rect 10870 22992 10876 23044
rect 10928 22992 10934 23044
rect 23842 23032 23848 23044
rect 23584 23004 23848 23032
rect 3145 22967 3203 22973
rect 3145 22933 3157 22967
rect 3191 22964 3203 22967
rect 4706 22964 4712 22976
rect 3191 22936 4712 22964
rect 3191 22933 3203 22936
rect 3145 22927 3203 22933
rect 4706 22924 4712 22936
rect 4764 22924 4770 22976
rect 12713 22967 12771 22973
rect 12713 22933 12725 22967
rect 12759 22964 12771 22967
rect 12986 22964 12992 22976
rect 12759 22936 12992 22964
rect 12759 22933 12771 22936
rect 12713 22927 12771 22933
rect 12986 22924 12992 22936
rect 13044 22924 13050 22976
rect 18782 22964 18788 22976
rect 18743 22936 18788 22964
rect 18782 22924 18788 22936
rect 18840 22924 18846 22976
rect 23385 22967 23443 22973
rect 23385 22933 23397 22967
rect 23431 22964 23443 22967
rect 23474 22964 23480 22976
rect 23431 22936 23480 22964
rect 23431 22933 23443 22936
rect 23385 22927 23443 22933
rect 23474 22924 23480 22936
rect 23532 22924 23538 22976
rect 23584 22973 23612 23004
rect 23842 22992 23848 23004
rect 23900 23032 23906 23044
rect 27798 23032 27804 23044
rect 23900 23004 27804 23032
rect 23900 22992 23906 23004
rect 27798 22992 27804 23004
rect 27856 22992 27862 23044
rect 28828 23032 28856 23063
rect 30926 23060 30932 23072
rect 30984 23060 30990 23112
rect 31018 23060 31024 23112
rect 31076 23100 31082 23112
rect 32401 23103 32459 23109
rect 32401 23100 32413 23103
rect 31076 23072 32413 23100
rect 31076 23060 31082 23072
rect 32401 23069 32413 23072
rect 32447 23100 32459 23103
rect 33321 23103 33379 23109
rect 33321 23100 33333 23103
rect 32447 23072 33333 23100
rect 32447 23069 32459 23072
rect 32401 23063 32459 23069
rect 33321 23069 33333 23072
rect 33367 23069 33379 23103
rect 33321 23063 33379 23069
rect 33413 23103 33471 23109
rect 33413 23069 33425 23103
rect 33459 23069 33471 23103
rect 33413 23063 33471 23069
rect 30006 23032 30012 23044
rect 28828 23004 30012 23032
rect 30006 22992 30012 23004
rect 30064 22992 30070 23044
rect 33428 23032 33456 23063
rect 33336 23004 33456 23032
rect 23569 22967 23627 22973
rect 23569 22933 23581 22967
rect 23615 22933 23627 22967
rect 23569 22927 23627 22933
rect 27522 22924 27528 22976
rect 27580 22964 27586 22976
rect 27617 22967 27675 22973
rect 27617 22964 27629 22967
rect 27580 22936 27629 22964
rect 27580 22924 27586 22936
rect 27617 22933 27629 22936
rect 27663 22933 27675 22967
rect 27617 22927 27675 22933
rect 28353 22967 28411 22973
rect 28353 22933 28365 22967
rect 28399 22964 28411 22967
rect 28534 22964 28540 22976
rect 28399 22936 28540 22964
rect 28399 22933 28411 22936
rect 28353 22927 28411 22933
rect 28534 22924 28540 22936
rect 28592 22924 28598 22976
rect 31386 22924 31392 22976
rect 31444 22964 31450 22976
rect 33336 22964 33364 23004
rect 31444 22936 33364 22964
rect 31444 22924 31450 22936
rect 1104 22874 34316 22896
rect 1104 22822 6517 22874
rect 6569 22822 6581 22874
rect 6633 22822 6645 22874
rect 6697 22822 6709 22874
rect 6761 22822 17588 22874
rect 17640 22822 17652 22874
rect 17704 22822 17716 22874
rect 17768 22822 17780 22874
rect 17832 22822 28658 22874
rect 28710 22822 28722 22874
rect 28774 22822 28786 22874
rect 28838 22822 28850 22874
rect 28902 22822 34316 22874
rect 1104 22800 34316 22822
rect 3326 22720 3332 22772
rect 3384 22760 3390 22772
rect 3421 22763 3479 22769
rect 3421 22760 3433 22763
rect 3384 22732 3433 22760
rect 3384 22720 3390 22732
rect 3421 22729 3433 22732
rect 3467 22729 3479 22763
rect 4154 22760 4160 22772
rect 4115 22732 4160 22760
rect 3421 22723 3479 22729
rect 4154 22720 4160 22732
rect 4212 22720 4218 22772
rect 6914 22760 6920 22772
rect 6875 22732 6920 22760
rect 6914 22720 6920 22732
rect 6972 22720 6978 22772
rect 10226 22720 10232 22772
rect 10284 22760 10290 22772
rect 10962 22760 10968 22772
rect 10284 22732 10968 22760
rect 10284 22720 10290 22732
rect 10962 22720 10968 22732
rect 11020 22720 11026 22772
rect 12986 22760 12992 22772
rect 12268 22732 12992 22760
rect 2682 22652 2688 22704
rect 2740 22692 2746 22704
rect 5810 22692 5816 22704
rect 2740 22664 5672 22692
rect 5771 22664 5816 22692
rect 2740 22652 2746 22664
rect 2700 22596 4476 22624
rect 2700 22568 2728 22596
rect 4448 22568 4476 22596
rect 4706 22584 4712 22636
rect 4764 22624 4770 22636
rect 4801 22627 4859 22633
rect 4801 22624 4813 22627
rect 4764 22596 4813 22624
rect 4764 22584 4770 22596
rect 4801 22593 4813 22596
rect 4847 22624 4859 22627
rect 5644 22624 5672 22664
rect 5810 22652 5816 22664
rect 5868 22652 5874 22704
rect 7006 22624 7012 22636
rect 4847 22596 5580 22624
rect 5644 22596 7012 22624
rect 4847 22593 4859 22596
rect 4801 22587 4859 22593
rect 2682 22556 2688 22568
rect 2595 22528 2688 22556
rect 2682 22516 2688 22528
rect 2740 22516 2746 22568
rect 2869 22559 2927 22565
rect 2869 22525 2881 22559
rect 2915 22556 2927 22559
rect 2958 22556 2964 22568
rect 2915 22528 2964 22556
rect 2915 22525 2927 22528
rect 2869 22519 2927 22525
rect 2958 22516 2964 22528
rect 3016 22516 3022 22568
rect 3326 22556 3332 22568
rect 3287 22528 3332 22556
rect 3326 22516 3332 22528
rect 3384 22516 3390 22568
rect 3513 22559 3571 22565
rect 3513 22525 3525 22559
rect 3559 22525 3571 22559
rect 4338 22556 4344 22568
rect 4299 22528 4344 22556
rect 3513 22519 3571 22525
rect 2774 22380 2780 22432
rect 2832 22420 2838 22432
rect 3528 22420 3556 22519
rect 4338 22516 4344 22528
rect 4396 22516 4402 22568
rect 4430 22516 4436 22568
rect 4488 22556 4494 22568
rect 5552 22565 5580 22596
rect 7006 22584 7012 22596
rect 7064 22624 7070 22636
rect 7926 22624 7932 22636
rect 7064 22596 7932 22624
rect 7064 22584 7070 22596
rect 5537 22559 5595 22565
rect 4488 22528 4533 22556
rect 4488 22516 4494 22528
rect 5537 22525 5549 22559
rect 5583 22525 5595 22559
rect 5537 22519 5595 22525
rect 5813 22559 5871 22565
rect 5813 22525 5825 22559
rect 5859 22556 5871 22559
rect 6270 22556 6276 22568
rect 5859 22528 6276 22556
rect 5859 22525 5871 22528
rect 5813 22519 5871 22525
rect 6270 22516 6276 22528
rect 6328 22516 6334 22568
rect 7300 22542 7328 22596
rect 7926 22584 7932 22596
rect 7984 22584 7990 22636
rect 8386 22624 8392 22636
rect 8347 22596 8392 22624
rect 8386 22584 8392 22596
rect 8444 22584 8450 22636
rect 8665 22627 8723 22633
rect 8665 22593 8677 22627
rect 8711 22624 8723 22627
rect 8754 22624 8760 22636
rect 8711 22596 8760 22624
rect 8711 22593 8723 22596
rect 8665 22587 8723 22593
rect 8754 22584 8760 22596
rect 8812 22584 8818 22636
rect 9125 22559 9183 22565
rect 9125 22525 9137 22559
rect 9171 22525 9183 22559
rect 9125 22519 9183 22525
rect 11057 22559 11115 22565
rect 11057 22525 11069 22559
rect 11103 22556 11115 22559
rect 11146 22556 11152 22568
rect 11103 22528 11152 22556
rect 11103 22525 11115 22528
rect 11057 22519 11115 22525
rect 4706 22488 4712 22500
rect 4667 22460 4712 22488
rect 4706 22448 4712 22460
rect 4764 22448 4770 22500
rect 9140 22488 9168 22519
rect 11146 22516 11152 22528
rect 11204 22556 11210 22568
rect 12268 22565 12296 22732
rect 12986 22720 12992 22732
rect 13044 22720 13050 22772
rect 15010 22720 15016 22772
rect 15068 22760 15074 22772
rect 15562 22760 15568 22772
rect 15068 22732 15568 22760
rect 15068 22720 15074 22732
rect 15562 22720 15568 22732
rect 15620 22760 15626 22772
rect 15841 22763 15899 22769
rect 15841 22760 15853 22763
rect 15620 22732 15853 22760
rect 15620 22720 15626 22732
rect 15841 22729 15853 22732
rect 15887 22729 15899 22763
rect 19518 22760 19524 22772
rect 19479 22732 19524 22760
rect 15841 22723 15899 22729
rect 19518 22720 19524 22732
rect 19576 22720 19582 22772
rect 26789 22763 26847 22769
rect 26789 22729 26801 22763
rect 26835 22760 26847 22763
rect 28258 22760 28264 22772
rect 26835 22732 28264 22760
rect 26835 22729 26847 22732
rect 26789 22723 26847 22729
rect 28258 22720 28264 22732
rect 28316 22720 28322 22772
rect 29822 22760 29828 22772
rect 28368 22732 29828 22760
rect 12526 22652 12532 22704
rect 12584 22692 12590 22704
rect 13081 22695 13139 22701
rect 13081 22692 13093 22695
rect 12584 22664 13093 22692
rect 12584 22652 12590 22664
rect 13081 22661 13093 22664
rect 13127 22661 13139 22695
rect 13081 22655 13139 22661
rect 19610 22652 19616 22704
rect 19668 22692 19674 22704
rect 21818 22692 21824 22704
rect 19668 22664 21824 22692
rect 19668 22652 19674 22664
rect 21818 22652 21824 22664
rect 21876 22652 21882 22704
rect 23566 22692 23572 22704
rect 22756 22664 23572 22692
rect 13170 22624 13176 22636
rect 13131 22596 13176 22624
rect 13170 22584 13176 22596
rect 13228 22584 13234 22636
rect 13814 22584 13820 22636
rect 13872 22624 13878 22636
rect 14093 22627 14151 22633
rect 14093 22624 14105 22627
rect 13872 22596 14105 22624
rect 13872 22584 13878 22596
rect 14093 22593 14105 22596
rect 14139 22624 14151 22627
rect 16298 22624 16304 22636
rect 14139 22596 16304 22624
rect 14139 22593 14151 22596
rect 14093 22587 14151 22593
rect 16298 22584 16304 22596
rect 16356 22584 16362 22636
rect 18782 22624 18788 22636
rect 18743 22596 18788 22624
rect 18782 22584 18788 22596
rect 18840 22584 18846 22636
rect 19705 22627 19763 22633
rect 19705 22593 19717 22627
rect 19751 22624 19763 22627
rect 20533 22627 20591 22633
rect 20533 22624 20545 22627
rect 19751 22596 20545 22624
rect 19751 22593 19763 22596
rect 19705 22587 19763 22593
rect 20533 22593 20545 22596
rect 20579 22624 20591 22627
rect 20579 22596 22094 22624
rect 20579 22593 20591 22596
rect 20533 22587 20591 22593
rect 12069 22559 12127 22565
rect 12069 22556 12081 22559
rect 11204 22528 12081 22556
rect 11204 22516 11210 22528
rect 12069 22525 12081 22528
rect 12115 22525 12127 22559
rect 12069 22519 12127 22525
rect 12253 22559 12311 22565
rect 12253 22525 12265 22559
rect 12299 22525 12311 22559
rect 12897 22559 12955 22565
rect 12897 22556 12909 22559
rect 12253 22519 12311 22525
rect 12406 22528 12909 22556
rect 8036 22460 9168 22488
rect 8036 22432 8064 22460
rect 10962 22448 10968 22500
rect 11020 22488 11026 22500
rect 12406 22488 12434 22528
rect 12897 22525 12909 22528
rect 12943 22556 12955 22559
rect 13354 22556 13360 22568
rect 12943 22528 13360 22556
rect 12943 22525 12955 22528
rect 12897 22519 12955 22525
rect 13354 22516 13360 22528
rect 13412 22516 13418 22568
rect 15470 22516 15476 22568
rect 15528 22516 15534 22568
rect 19061 22559 19119 22565
rect 19061 22525 19073 22559
rect 19107 22556 19119 22559
rect 19426 22556 19432 22568
rect 19107 22528 19432 22556
rect 19107 22525 19119 22528
rect 19061 22519 19119 22525
rect 19426 22516 19432 22528
rect 19484 22516 19490 22568
rect 19521 22559 19579 22565
rect 19521 22525 19533 22559
rect 19567 22525 19579 22559
rect 19521 22519 19579 22525
rect 19889 22559 19947 22565
rect 19889 22525 19901 22559
rect 19935 22556 19947 22559
rect 19978 22556 19984 22568
rect 19935 22528 19984 22556
rect 19935 22525 19947 22528
rect 19889 22519 19947 22525
rect 14366 22488 14372 22500
rect 11020 22460 12434 22488
rect 14327 22460 14372 22488
rect 11020 22448 11026 22460
rect 14366 22448 14372 22460
rect 14424 22448 14430 22500
rect 19334 22488 19340 22500
rect 18354 22460 19340 22488
rect 19334 22448 19340 22460
rect 19392 22448 19398 22500
rect 6730 22420 6736 22432
rect 2832 22392 2877 22420
rect 3528 22392 6736 22420
rect 2832 22380 2838 22392
rect 6730 22380 6736 22392
rect 6788 22380 6794 22432
rect 8018 22380 8024 22432
rect 8076 22380 8082 22432
rect 9306 22420 9312 22432
rect 9267 22392 9312 22420
rect 9306 22380 9312 22392
rect 9364 22380 9370 22432
rect 11790 22380 11796 22432
rect 11848 22420 11854 22432
rect 12161 22423 12219 22429
rect 12161 22420 12173 22423
rect 11848 22392 12173 22420
rect 11848 22380 11854 22392
rect 12161 22389 12173 22392
rect 12207 22389 12219 22423
rect 17310 22420 17316 22432
rect 17223 22392 17316 22420
rect 12161 22383 12219 22389
rect 17310 22380 17316 22392
rect 17368 22420 17374 22432
rect 19536 22420 19564 22519
rect 19978 22516 19984 22528
rect 20036 22556 20042 22568
rect 20349 22559 20407 22565
rect 20349 22556 20361 22559
rect 20036 22528 20361 22556
rect 20036 22516 20042 22528
rect 20349 22525 20361 22528
rect 20395 22525 20407 22559
rect 20717 22559 20775 22565
rect 20717 22556 20729 22559
rect 20349 22519 20407 22525
rect 20548 22528 20729 22556
rect 20548 22500 20576 22528
rect 20717 22525 20729 22528
rect 20763 22525 20775 22559
rect 20717 22519 20775 22525
rect 19702 22448 19708 22500
rect 19760 22488 19766 22500
rect 20530 22488 20536 22500
rect 19760 22460 20536 22488
rect 19760 22448 19766 22460
rect 20530 22448 20536 22460
rect 20588 22448 20594 22500
rect 22066 22488 22094 22596
rect 22756 22565 22784 22664
rect 23566 22652 23572 22664
rect 23624 22652 23630 22704
rect 23753 22695 23811 22701
rect 23753 22661 23765 22695
rect 23799 22661 23811 22695
rect 28368 22692 28396 22732
rect 29822 22720 29828 22732
rect 29880 22720 29886 22772
rect 30006 22760 30012 22772
rect 29967 22732 30012 22760
rect 30006 22720 30012 22732
rect 30064 22720 30070 22772
rect 30837 22763 30895 22769
rect 30837 22729 30849 22763
rect 30883 22760 30895 22763
rect 30926 22760 30932 22772
rect 30883 22732 30932 22760
rect 30883 22729 30895 22732
rect 30837 22723 30895 22729
rect 30926 22720 30932 22732
rect 30984 22720 30990 22772
rect 23753 22655 23811 22661
rect 25792 22664 28396 22692
rect 23768 22624 23796 22655
rect 24673 22627 24731 22633
rect 24673 22624 24685 22627
rect 23768 22596 24685 22624
rect 24673 22593 24685 22596
rect 24719 22593 24731 22627
rect 24673 22587 24731 22593
rect 24762 22584 24768 22636
rect 24820 22624 24826 22636
rect 25792 22624 25820 22664
rect 27062 22624 27068 22636
rect 24820 22596 25820 22624
rect 24820 22584 24826 22596
rect 22741 22559 22799 22565
rect 22741 22525 22753 22559
rect 22787 22525 22799 22559
rect 22741 22519 22799 22525
rect 22925 22559 22983 22565
rect 22925 22525 22937 22559
rect 22971 22525 22983 22559
rect 22925 22519 22983 22525
rect 22833 22491 22891 22497
rect 22833 22488 22845 22491
rect 22066 22460 22845 22488
rect 22833 22457 22845 22460
rect 22879 22457 22891 22491
rect 22833 22451 22891 22457
rect 17368 22392 19564 22420
rect 19797 22423 19855 22429
rect 17368 22380 17374 22392
rect 19797 22389 19809 22423
rect 19843 22420 19855 22423
rect 19886 22420 19892 22432
rect 19843 22392 19892 22420
rect 19843 22389 19855 22392
rect 19797 22383 19855 22389
rect 19886 22380 19892 22392
rect 19944 22420 19950 22432
rect 20346 22420 20352 22432
rect 19944 22392 20352 22420
rect 19944 22380 19950 22392
rect 20346 22380 20352 22392
rect 20404 22420 20410 22432
rect 20441 22423 20499 22429
rect 20441 22420 20453 22423
rect 20404 22392 20453 22420
rect 20404 22380 20410 22392
rect 20441 22389 20453 22392
rect 20487 22389 20499 22423
rect 20622 22420 20628 22432
rect 20583 22392 20628 22420
rect 20441 22383 20499 22389
rect 20622 22380 20628 22392
rect 20680 22380 20686 22432
rect 22940 22420 22968 22519
rect 23014 22516 23020 22568
rect 23072 22556 23078 22568
rect 23385 22559 23443 22565
rect 23385 22556 23397 22559
rect 23072 22528 23397 22556
rect 23072 22516 23078 22528
rect 23385 22525 23397 22528
rect 23431 22525 23443 22559
rect 23385 22519 23443 22525
rect 23477 22559 23535 22565
rect 23477 22525 23489 22559
rect 23523 22556 23535 22559
rect 23658 22556 23664 22568
rect 23523 22528 23664 22556
rect 23523 22525 23535 22528
rect 23477 22519 23535 22525
rect 23658 22516 23664 22528
rect 23716 22516 23722 22568
rect 23842 22556 23848 22568
rect 23803 22528 23848 22556
rect 23842 22516 23848 22528
rect 23900 22516 23906 22568
rect 23937 22559 23995 22565
rect 23937 22525 23949 22559
rect 23983 22556 23995 22559
rect 24026 22556 24032 22568
rect 23983 22528 24032 22556
rect 23983 22525 23995 22528
rect 23937 22519 23995 22525
rect 24026 22516 24032 22528
rect 24084 22516 24090 22568
rect 24394 22556 24400 22568
rect 24355 22528 24400 22556
rect 24394 22516 24400 22528
rect 24452 22516 24458 22568
rect 25792 22542 25820 22596
rect 26712 22596 27068 22624
rect 26712 22565 26740 22596
rect 27062 22584 27068 22596
rect 27120 22624 27126 22636
rect 27522 22624 27528 22636
rect 27120 22596 27528 22624
rect 27120 22584 27126 22596
rect 27522 22584 27528 22596
rect 27580 22584 27586 22636
rect 28534 22624 28540 22636
rect 28495 22596 28540 22624
rect 28534 22584 28540 22596
rect 28592 22584 28598 22636
rect 30024 22624 30052 22720
rect 30834 22624 30840 22636
rect 30024 22596 30840 22624
rect 30834 22584 30840 22596
rect 30892 22624 30898 22636
rect 31386 22624 31392 22636
rect 30892 22596 31248 22624
rect 31347 22596 31392 22624
rect 30892 22584 30898 22596
rect 26697 22559 26755 22565
rect 26697 22525 26709 22559
rect 26743 22525 26755 22559
rect 26697 22519 26755 22525
rect 26878 22516 26884 22568
rect 26936 22556 26942 22568
rect 28261 22559 28319 22565
rect 28261 22556 28273 22559
rect 26936 22528 28273 22556
rect 26936 22516 26942 22528
rect 28261 22525 28273 22528
rect 28307 22525 28319 22559
rect 31220 22556 31248 22596
rect 31386 22584 31392 22596
rect 31444 22584 31450 22636
rect 31297 22559 31355 22565
rect 31297 22556 31309 22559
rect 31220 22528 31309 22556
rect 28261 22519 28319 22525
rect 31297 22525 31309 22528
rect 31343 22525 31355 22559
rect 31297 22519 31355 22525
rect 23934 22420 23940 22432
rect 22940 22392 23940 22420
rect 23934 22380 23940 22392
rect 23992 22380 23998 22432
rect 26142 22420 26148 22432
rect 26103 22392 26148 22420
rect 26142 22380 26148 22392
rect 26200 22380 26206 22432
rect 28276 22420 28304 22519
rect 29822 22488 29828 22500
rect 29735 22460 29828 22488
rect 29822 22448 29828 22460
rect 29880 22488 29886 22500
rect 32582 22488 32588 22500
rect 29880 22460 32588 22488
rect 29880 22448 29886 22460
rect 32582 22448 32588 22460
rect 32640 22448 32646 22500
rect 29362 22420 29368 22432
rect 28276 22392 29368 22420
rect 29362 22380 29368 22392
rect 29420 22380 29426 22432
rect 30926 22380 30932 22432
rect 30984 22420 30990 22432
rect 31205 22423 31263 22429
rect 31205 22420 31217 22423
rect 30984 22392 31217 22420
rect 30984 22380 30990 22392
rect 31205 22389 31217 22392
rect 31251 22389 31263 22423
rect 31205 22383 31263 22389
rect 1104 22330 34316 22352
rect 1104 22278 12052 22330
rect 12104 22278 12116 22330
rect 12168 22278 12180 22330
rect 12232 22278 12244 22330
rect 12296 22278 23123 22330
rect 23175 22278 23187 22330
rect 23239 22278 23251 22330
rect 23303 22278 23315 22330
rect 23367 22278 34316 22330
rect 1104 22256 34316 22278
rect 4706 22176 4712 22228
rect 4764 22216 4770 22228
rect 4801 22219 4859 22225
rect 4801 22216 4813 22219
rect 4764 22188 4813 22216
rect 4764 22176 4770 22188
rect 4801 22185 4813 22188
rect 4847 22185 4859 22219
rect 4801 22179 4859 22185
rect 10318 22176 10324 22228
rect 10376 22216 10382 22228
rect 10870 22216 10876 22228
rect 10376 22188 10876 22216
rect 10376 22176 10382 22188
rect 10870 22176 10876 22188
rect 10928 22216 10934 22228
rect 10965 22219 11023 22225
rect 10965 22216 10977 22219
rect 10928 22188 10977 22216
rect 10928 22176 10934 22188
rect 10965 22185 10977 22188
rect 11011 22216 11023 22219
rect 11698 22216 11704 22228
rect 11011 22188 11704 22216
rect 11011 22185 11023 22188
rect 10965 22179 11023 22185
rect 11698 22176 11704 22188
rect 11756 22176 11762 22228
rect 12342 22216 12348 22228
rect 12303 22188 12348 22216
rect 12342 22176 12348 22188
rect 12400 22176 12406 22228
rect 16574 22176 16580 22228
rect 16632 22176 16638 22228
rect 21450 22176 21456 22228
rect 21508 22216 21514 22228
rect 21508 22188 21680 22216
rect 21508 22176 21514 22188
rect 2682 22108 2688 22160
rect 2740 22148 2746 22160
rect 2740 22120 3004 22148
rect 2740 22108 2746 22120
rect 2976 22089 3004 22120
rect 3326 22108 3332 22160
rect 3384 22148 3390 22160
rect 4246 22148 4252 22160
rect 3384 22120 4252 22148
rect 3384 22108 3390 22120
rect 4246 22108 4252 22120
rect 4304 22148 4310 22160
rect 4304 22120 6500 22148
rect 4304 22108 4310 22120
rect 2961 22083 3019 22089
rect 2961 22049 2973 22083
rect 3007 22049 3019 22083
rect 2961 22043 3019 22049
rect 4614 22040 4620 22092
rect 4672 22080 4678 22092
rect 4709 22083 4767 22089
rect 4709 22080 4721 22083
rect 4672 22052 4721 22080
rect 4672 22040 4678 22052
rect 4709 22049 4721 22052
rect 4755 22049 4767 22083
rect 4890 22080 4896 22092
rect 4851 22052 4896 22080
rect 4709 22043 4767 22049
rect 4890 22040 4896 22052
rect 4948 22040 4954 22092
rect 5350 22080 5356 22092
rect 5311 22052 5356 22080
rect 5350 22040 5356 22052
rect 5408 22040 5414 22092
rect 5534 22080 5540 22092
rect 5495 22052 5540 22080
rect 5534 22040 5540 22052
rect 5592 22040 5598 22092
rect 6472 22089 6500 22120
rect 6730 22108 6736 22160
rect 6788 22148 6794 22160
rect 6788 22120 7236 22148
rect 6788 22108 6794 22120
rect 6457 22083 6515 22089
rect 6457 22049 6469 22083
rect 6503 22049 6515 22083
rect 6914 22080 6920 22092
rect 6875 22052 6920 22080
rect 6457 22043 6515 22049
rect 6914 22040 6920 22052
rect 6972 22040 6978 22092
rect 7208 22089 7236 22120
rect 9306 22108 9312 22160
rect 9364 22148 9370 22160
rect 11054 22148 11060 22160
rect 9364 22120 11060 22148
rect 9364 22108 9370 22120
rect 11054 22108 11060 22120
rect 11112 22148 11118 22160
rect 13814 22148 13820 22160
rect 11112 22120 13820 22148
rect 11112 22108 11118 22120
rect 13814 22108 13820 22120
rect 13872 22108 13878 22160
rect 16592 22148 16620 22176
rect 16408 22120 16620 22148
rect 16669 22151 16727 22157
rect 7193 22083 7251 22089
rect 7193 22049 7205 22083
rect 7239 22080 7251 22083
rect 7466 22080 7472 22092
rect 7239 22052 7472 22080
rect 7239 22049 7251 22052
rect 7193 22043 7251 22049
rect 7466 22040 7472 22052
rect 7524 22040 7530 22092
rect 7926 22040 7932 22092
rect 7984 22080 7990 22092
rect 10778 22080 10784 22092
rect 7984 22052 10784 22080
rect 7984 22040 7990 22052
rect 10778 22040 10784 22052
rect 10836 22040 10842 22092
rect 11146 22080 11152 22092
rect 11107 22052 11152 22080
rect 11146 22040 11152 22052
rect 11204 22040 11210 22092
rect 12342 22080 12348 22092
rect 12303 22052 12348 22080
rect 12342 22040 12348 22052
rect 12400 22040 12406 22092
rect 13354 22080 13360 22092
rect 13315 22052 13360 22080
rect 13354 22040 13360 22052
rect 13412 22040 13418 22092
rect 15286 22080 15292 22092
rect 13648 22052 15292 22080
rect 2685 22015 2743 22021
rect 2685 21981 2697 22015
rect 2731 22012 2743 22015
rect 2774 22012 2780 22024
rect 2731 21984 2780 22012
rect 2731 21981 2743 21984
rect 2685 21975 2743 21981
rect 2774 21972 2780 21984
rect 2832 21972 2838 22024
rect 4062 21972 4068 22024
rect 4120 22012 4126 22024
rect 5368 22012 5396 22040
rect 7098 22012 7104 22024
rect 4120 21984 5396 22012
rect 7059 21984 7104 22012
rect 4120 21972 4126 21984
rect 7098 21972 7104 21984
rect 7156 21972 7162 22024
rect 11882 21972 11888 22024
rect 11940 22012 11946 22024
rect 11977 22015 12035 22021
rect 11977 22012 11989 22015
rect 11940 21984 11989 22012
rect 11940 21972 11946 21984
rect 11977 21981 11989 21984
rect 12023 21981 12035 22015
rect 12526 22012 12532 22024
rect 12487 21984 12532 22012
rect 11977 21975 12035 21981
rect 12526 21972 12532 21984
rect 12584 21972 12590 22024
rect 13648 22021 13676 22052
rect 15286 22040 15292 22052
rect 15344 22040 15350 22092
rect 16408 22089 16436 22120
rect 16669 22117 16681 22151
rect 16715 22148 16727 22151
rect 18598 22148 18604 22160
rect 16715 22120 18604 22148
rect 16715 22117 16727 22120
rect 16669 22111 16727 22117
rect 18598 22108 18604 22120
rect 18656 22108 18662 22160
rect 21652 22148 21680 22188
rect 30668 22188 31754 22216
rect 21726 22148 21732 22160
rect 21652 22134 21732 22148
rect 21666 22120 21732 22134
rect 21726 22108 21732 22120
rect 21784 22108 21790 22160
rect 21818 22108 21824 22160
rect 21876 22148 21882 22160
rect 22361 22151 22419 22157
rect 22361 22148 22373 22151
rect 21876 22120 22373 22148
rect 21876 22108 21882 22120
rect 22361 22117 22373 22120
rect 22407 22117 22419 22151
rect 22361 22111 22419 22117
rect 22756 22120 24808 22148
rect 22756 22092 22784 22120
rect 16393 22083 16451 22089
rect 16393 22049 16405 22083
rect 16439 22080 16451 22083
rect 16574 22080 16580 22092
rect 16439 22052 16473 22080
rect 16535 22052 16580 22080
rect 16439 22049 16451 22052
rect 16393 22043 16451 22049
rect 16574 22040 16580 22052
rect 16632 22040 16638 22092
rect 22738 22080 22744 22092
rect 22651 22052 22744 22080
rect 22738 22040 22744 22052
rect 22796 22040 22802 22092
rect 23385 22083 23443 22089
rect 23385 22049 23397 22083
rect 23431 22080 23443 22083
rect 23566 22080 23572 22092
rect 23431 22052 23572 22080
rect 23431 22049 23443 22052
rect 23385 22043 23443 22049
rect 23566 22040 23572 22052
rect 23624 22080 23630 22092
rect 24394 22080 24400 22092
rect 23624 22052 24400 22080
rect 23624 22040 23630 22052
rect 24394 22040 24400 22052
rect 24452 22040 24458 22092
rect 24780 22024 24808 22120
rect 27632 22120 27844 22148
rect 25774 22040 25780 22092
rect 25832 22080 25838 22092
rect 25961 22083 26019 22089
rect 25961 22080 25973 22083
rect 25832 22052 25973 22080
rect 25832 22040 25838 22052
rect 25961 22049 25973 22052
rect 26007 22049 26019 22083
rect 25961 22043 26019 22049
rect 26142 22040 26148 22092
rect 26200 22080 26206 22092
rect 26421 22083 26479 22089
rect 26421 22080 26433 22083
rect 26200 22052 26433 22080
rect 26200 22040 26206 22052
rect 26421 22049 26433 22052
rect 26467 22049 26479 22083
rect 27062 22080 27068 22092
rect 26421 22043 26479 22049
rect 26528 22052 26832 22080
rect 27023 22052 27068 22080
rect 13633 22015 13691 22021
rect 13633 21981 13645 22015
rect 13679 21981 13691 22015
rect 13633 21975 13691 21981
rect 19426 21972 19432 22024
rect 19484 22012 19490 22024
rect 20162 22012 20168 22024
rect 19484 21984 20168 22012
rect 19484 21972 19490 21984
rect 20162 21972 20168 21984
rect 20220 21972 20226 22024
rect 20441 22015 20499 22021
rect 20441 21981 20453 22015
rect 20487 22012 20499 22015
rect 22370 22012 22376 22024
rect 20487 21984 22376 22012
rect 20487 21981 20499 21984
rect 20441 21975 20499 21981
rect 22370 21972 22376 21984
rect 22428 21972 22434 22024
rect 23753 22015 23811 22021
rect 7282 21904 7288 21956
rect 7340 21944 7346 21956
rect 12158 21944 12164 21956
rect 7340 21916 12164 21944
rect 7340 21904 7346 21916
rect 12158 21904 12164 21916
rect 12216 21904 12222 21956
rect 13449 21947 13507 21953
rect 13449 21944 13461 21947
rect 12406 21916 13461 21944
rect 1670 21836 1676 21888
rect 1728 21876 1734 21888
rect 2777 21879 2835 21885
rect 2777 21876 2789 21879
rect 1728 21848 2789 21876
rect 1728 21836 1734 21848
rect 2777 21845 2789 21848
rect 2823 21845 2835 21879
rect 2777 21839 2835 21845
rect 2869 21879 2927 21885
rect 2869 21845 2881 21879
rect 2915 21876 2927 21879
rect 2958 21876 2964 21888
rect 2915 21848 2964 21876
rect 2915 21845 2927 21848
rect 2869 21839 2927 21845
rect 2958 21836 2964 21848
rect 3016 21836 3022 21888
rect 4982 21836 4988 21888
rect 5040 21876 5046 21888
rect 5537 21879 5595 21885
rect 5537 21876 5549 21879
rect 5040 21848 5549 21876
rect 5040 21836 5046 21848
rect 5537 21845 5549 21848
rect 5583 21845 5595 21879
rect 5537 21839 5595 21845
rect 11238 21836 11244 21888
rect 11296 21876 11302 21888
rect 12406 21876 12434 21916
rect 13449 21913 13461 21916
rect 13495 21913 13507 21947
rect 13449 21907 13507 21913
rect 21818 21904 21824 21956
rect 21876 21944 21882 21956
rect 23032 21944 23060 21998
rect 23753 21981 23765 22015
rect 23799 22012 23811 22015
rect 23934 22012 23940 22024
rect 23799 21984 23940 22012
rect 23799 21981 23811 21984
rect 23753 21975 23811 21981
rect 23934 21972 23940 21984
rect 23992 22012 23998 22024
rect 24486 22012 24492 22024
rect 23992 21984 24492 22012
rect 23992 21972 23998 21984
rect 24486 21972 24492 21984
rect 24544 21972 24550 22024
rect 24762 21972 24768 22024
rect 24820 22012 24826 22024
rect 26528 22012 26556 22052
rect 24820 21984 26556 22012
rect 26697 22015 26755 22021
rect 24820 21972 24826 21984
rect 26697 21981 26709 22015
rect 26743 21981 26755 22015
rect 26697 21975 26755 21981
rect 26712 21944 26740 21975
rect 21876 21916 26740 21944
rect 26804 21944 26832 22052
rect 27062 22040 27068 22052
rect 27120 22040 27126 22092
rect 27430 22080 27436 22092
rect 27343 22052 27436 22080
rect 27430 22040 27436 22052
rect 27488 22080 27494 22092
rect 27632 22080 27660 22120
rect 27488 22052 27660 22080
rect 27709 22083 27767 22089
rect 27488 22040 27494 22052
rect 27709 22049 27721 22083
rect 27755 22049 27767 22083
rect 27816 22080 27844 22120
rect 28166 22108 28172 22160
rect 28224 22148 28230 22160
rect 30668 22157 30696 22188
rect 30653 22151 30711 22157
rect 28224 22120 28672 22148
rect 28224 22108 28230 22120
rect 28644 22089 28672 22120
rect 30653 22117 30665 22151
rect 30699 22117 30711 22151
rect 30653 22111 30711 22117
rect 30834 22108 30840 22160
rect 30892 22157 30898 22160
rect 30892 22151 30916 22157
rect 30904 22117 30916 22151
rect 31726 22148 31754 22188
rect 31846 22148 31852 22160
rect 31726 22120 31852 22148
rect 30892 22111 30916 22117
rect 30892 22108 30898 22111
rect 31846 22108 31852 22120
rect 31904 22108 31910 22160
rect 28261 22083 28319 22089
rect 28261 22080 28273 22083
rect 27816 22052 28273 22080
rect 27709 22043 27767 22049
rect 28261 22049 28273 22052
rect 28307 22049 28319 22083
rect 28261 22043 28319 22049
rect 28629 22083 28687 22089
rect 28629 22049 28641 22083
rect 28675 22049 28687 22083
rect 28629 22043 28687 22049
rect 29273 22083 29331 22089
rect 29273 22049 29285 22083
rect 29319 22049 29331 22083
rect 29273 22043 29331 22049
rect 31665 22083 31723 22089
rect 31665 22049 31677 22083
rect 31711 22049 31723 22083
rect 32030 22080 32036 22092
rect 31991 22052 32036 22080
rect 31665 22043 31723 22049
rect 27724 22012 27752 22043
rect 27982 22012 27988 22024
rect 27724 21984 27988 22012
rect 27982 21972 27988 21984
rect 28040 22012 28046 22024
rect 29288 22012 29316 22043
rect 31481 22015 31539 22021
rect 31481 22012 31493 22015
rect 28040 21984 31493 22012
rect 28040 21972 28046 21984
rect 31481 21981 31493 21984
rect 31527 21981 31539 22015
rect 31481 21975 31539 21981
rect 30650 21944 30656 21956
rect 26804 21916 30656 21944
rect 21876 21904 21882 21916
rect 30650 21904 30656 21916
rect 30708 21904 30714 21956
rect 31021 21947 31079 21953
rect 31021 21913 31033 21947
rect 31067 21944 31079 21947
rect 31680 21944 31708 22043
rect 32030 22040 32036 22052
rect 32088 22040 32094 22092
rect 32677 22083 32735 22089
rect 32677 22049 32689 22083
rect 32723 22080 32735 22083
rect 33042 22080 33048 22092
rect 32723 22052 33048 22080
rect 32723 22049 32735 22052
rect 32677 22043 32735 22049
rect 33042 22040 33048 22052
rect 33100 22040 33106 22092
rect 31067 21916 31708 21944
rect 31067 21913 31079 21916
rect 31021 21907 31079 21913
rect 11296 21848 12434 21876
rect 13541 21879 13599 21885
rect 11296 21836 11302 21848
rect 13541 21845 13553 21879
rect 13587 21876 13599 21879
rect 14826 21876 14832 21888
rect 13587 21848 14832 21876
rect 13587 21845 13599 21848
rect 13541 21839 13599 21845
rect 14826 21836 14832 21848
rect 14884 21836 14890 21888
rect 21910 21876 21916 21888
rect 21871 21848 21916 21876
rect 21910 21836 21916 21848
rect 21968 21836 21974 21888
rect 26510 21836 26516 21888
rect 26568 21876 26574 21888
rect 28353 21879 28411 21885
rect 28353 21876 28365 21879
rect 26568 21848 28365 21876
rect 26568 21836 26574 21848
rect 28353 21845 28365 21848
rect 28399 21876 28411 21879
rect 29638 21876 29644 21888
rect 28399 21848 29644 21876
rect 28399 21845 28411 21848
rect 28353 21839 28411 21845
rect 29638 21836 29644 21848
rect 29696 21836 29702 21888
rect 30837 21879 30895 21885
rect 30837 21845 30849 21879
rect 30883 21876 30895 21879
rect 30926 21876 30932 21888
rect 30883 21848 30932 21876
rect 30883 21845 30895 21848
rect 30837 21839 30895 21845
rect 30926 21836 30932 21848
rect 30984 21836 30990 21888
rect 1104 21786 34316 21808
rect 1104 21734 6517 21786
rect 6569 21734 6581 21786
rect 6633 21734 6645 21786
rect 6697 21734 6709 21786
rect 6761 21734 17588 21786
rect 17640 21734 17652 21786
rect 17704 21734 17716 21786
rect 17768 21734 17780 21786
rect 17832 21734 28658 21786
rect 28710 21734 28722 21786
rect 28774 21734 28786 21786
rect 28838 21734 28850 21786
rect 28902 21734 34316 21786
rect 1104 21712 34316 21734
rect 11146 21672 11152 21684
rect 11107 21644 11152 21672
rect 11146 21632 11152 21644
rect 11204 21632 11210 21684
rect 12434 21632 12440 21684
rect 12492 21672 12498 21684
rect 12805 21675 12863 21681
rect 12805 21672 12817 21675
rect 12492 21644 12817 21672
rect 12492 21632 12498 21644
rect 12805 21641 12817 21644
rect 12851 21641 12863 21675
rect 19978 21672 19984 21684
rect 19939 21644 19984 21672
rect 12805 21635 12863 21641
rect 19978 21632 19984 21644
rect 20036 21632 20042 21684
rect 20714 21632 20720 21684
rect 20772 21672 20778 21684
rect 21269 21675 21327 21681
rect 21269 21672 21281 21675
rect 20772 21644 21281 21672
rect 20772 21632 20778 21644
rect 21269 21641 21281 21644
rect 21315 21641 21327 21675
rect 21269 21635 21327 21641
rect 21637 21675 21695 21681
rect 21637 21641 21649 21675
rect 21683 21672 21695 21675
rect 21910 21672 21916 21684
rect 21683 21644 21916 21672
rect 21683 21641 21695 21644
rect 21637 21635 21695 21641
rect 21910 21632 21916 21644
rect 21968 21632 21974 21684
rect 22370 21632 22376 21684
rect 22428 21672 22434 21684
rect 23201 21675 23259 21681
rect 23201 21672 23213 21675
rect 22428 21644 23213 21672
rect 22428 21632 22434 21644
rect 23201 21641 23213 21644
rect 23247 21641 23259 21675
rect 23201 21635 23259 21641
rect 23842 21632 23848 21684
rect 23900 21672 23906 21684
rect 24397 21675 24455 21681
rect 24397 21672 24409 21675
rect 23900 21644 24409 21672
rect 23900 21632 23906 21644
rect 24397 21641 24409 21644
rect 24443 21641 24455 21675
rect 24397 21635 24455 21641
rect 24486 21632 24492 21684
rect 24544 21672 24550 21684
rect 25317 21675 25375 21681
rect 25317 21672 25329 21675
rect 24544 21644 25329 21672
rect 24544 21632 24550 21644
rect 25317 21641 25329 21644
rect 25363 21641 25375 21675
rect 25498 21672 25504 21684
rect 25459 21644 25504 21672
rect 25317 21635 25375 21641
rect 25498 21632 25504 21644
rect 25556 21632 25562 21684
rect 29454 21672 29460 21684
rect 25608 21644 29460 21672
rect 11698 21564 11704 21616
rect 11756 21604 11762 21616
rect 11756 21576 12480 21604
rect 11756 21564 11762 21576
rect 1670 21536 1676 21548
rect 1631 21508 1676 21536
rect 1670 21496 1676 21508
rect 1728 21496 1734 21548
rect 3145 21539 3203 21545
rect 3145 21505 3157 21539
rect 3191 21536 3203 21539
rect 4154 21536 4160 21548
rect 3191 21508 4160 21536
rect 3191 21505 3203 21508
rect 3145 21499 3203 21505
rect 4154 21496 4160 21508
rect 4212 21496 4218 21548
rect 4798 21536 4804 21548
rect 4759 21508 4804 21536
rect 4798 21496 4804 21508
rect 4856 21496 4862 21548
rect 4982 21536 4988 21548
rect 4943 21508 4988 21536
rect 4982 21496 4988 21508
rect 5040 21496 5046 21548
rect 8849 21539 8907 21545
rect 8849 21505 8861 21539
rect 8895 21536 8907 21539
rect 10134 21536 10140 21548
rect 8895 21508 10140 21536
rect 8895 21505 8907 21508
rect 8849 21499 8907 21505
rect 10134 21496 10140 21508
rect 10192 21536 10198 21548
rect 11238 21536 11244 21548
rect 10192 21508 11244 21536
rect 10192 21496 10198 21508
rect 11238 21496 11244 21508
rect 11296 21496 11302 21548
rect 1394 21468 1400 21480
rect 1355 21440 1400 21468
rect 1394 21428 1400 21440
rect 1452 21428 1458 21480
rect 3050 21428 3056 21480
rect 3108 21468 3114 21480
rect 3878 21468 3884 21480
rect 3108 21440 3884 21468
rect 3108 21428 3114 21440
rect 3878 21428 3884 21440
rect 3936 21428 3942 21480
rect 4062 21468 4068 21480
rect 4023 21440 4068 21468
rect 4062 21428 4068 21440
rect 4120 21428 4126 21480
rect 8018 21468 8024 21480
rect 7979 21440 8024 21468
rect 8018 21428 8024 21440
rect 8076 21428 8082 21480
rect 8481 21471 8539 21477
rect 8481 21437 8493 21471
rect 8527 21437 8539 21471
rect 8662 21468 8668 21480
rect 8623 21440 8668 21468
rect 8481 21431 8539 21437
rect 2608 21344 2636 21386
rect 2590 21292 2596 21344
rect 2648 21292 2654 21344
rect 3970 21332 3976 21344
rect 3883 21304 3976 21332
rect 3970 21292 3976 21304
rect 4028 21332 4034 21344
rect 5077 21335 5135 21341
rect 5077 21332 5089 21335
rect 4028 21304 5089 21332
rect 4028 21292 4034 21304
rect 5077 21301 5089 21304
rect 5123 21301 5135 21335
rect 5077 21295 5135 21301
rect 5445 21335 5503 21341
rect 5445 21301 5457 21335
rect 5491 21332 5503 21335
rect 5718 21332 5724 21344
rect 5491 21304 5724 21332
rect 5491 21301 5503 21304
rect 5445 21295 5503 21301
rect 5718 21292 5724 21304
rect 5776 21292 5782 21344
rect 8202 21292 8208 21344
rect 8260 21332 8266 21344
rect 8496 21332 8524 21431
rect 8662 21428 8668 21440
rect 8720 21428 8726 21480
rect 8754 21428 8760 21480
rect 8812 21468 8818 21480
rect 9398 21468 9404 21480
rect 8812 21440 9404 21468
rect 8812 21428 8818 21440
rect 9398 21428 9404 21440
rect 9456 21428 9462 21480
rect 10778 21428 10784 21480
rect 10836 21428 10842 21480
rect 11790 21428 11796 21480
rect 11848 21468 11854 21480
rect 12452 21477 12480 21576
rect 12526 21564 12532 21616
rect 12584 21604 12590 21616
rect 24762 21604 24768 21616
rect 12584 21576 12664 21604
rect 24723 21576 24768 21604
rect 12584 21564 12590 21576
rect 12069 21471 12127 21477
rect 12069 21468 12081 21471
rect 11848 21440 12081 21468
rect 11848 21428 11854 21440
rect 12069 21437 12081 21440
rect 12115 21437 12127 21471
rect 12069 21431 12127 21437
rect 12257 21471 12315 21477
rect 12257 21437 12269 21471
rect 12303 21437 12315 21471
rect 12257 21431 12315 21437
rect 12348 21471 12406 21477
rect 12348 21437 12360 21471
rect 12394 21437 12406 21471
rect 12348 21431 12406 21437
rect 12437 21471 12495 21477
rect 12437 21437 12449 21471
rect 12483 21468 12495 21471
rect 12526 21468 12532 21480
rect 12483 21440 12532 21468
rect 12483 21437 12495 21440
rect 12437 21431 12495 21437
rect 9674 21400 9680 21412
rect 9635 21372 9680 21400
rect 9674 21360 9680 21372
rect 9732 21360 9738 21412
rect 12268 21400 12296 21431
rect 12366 21400 12394 21431
rect 12526 21428 12532 21440
rect 12584 21428 12590 21480
rect 12636 21477 12664 21576
rect 24762 21564 24768 21576
rect 24820 21564 24826 21616
rect 14366 21536 14372 21548
rect 14327 21508 14372 21536
rect 14366 21496 14372 21508
rect 14424 21496 14430 21548
rect 14734 21536 14740 21548
rect 14476 21508 14740 21536
rect 12621 21471 12679 21477
rect 12621 21437 12633 21471
rect 12667 21468 12679 21471
rect 12894 21468 12900 21480
rect 12667 21440 12900 21468
rect 12667 21437 12679 21440
rect 12621 21431 12679 21437
rect 12894 21428 12900 21440
rect 12952 21428 12958 21480
rect 13814 21468 13820 21480
rect 13775 21440 13820 21468
rect 13814 21428 13820 21440
rect 13872 21428 13878 21480
rect 14476 21477 14504 21508
rect 14734 21496 14740 21508
rect 14792 21496 14798 21548
rect 17773 21539 17831 21545
rect 17773 21505 17785 21539
rect 17819 21536 17831 21539
rect 19702 21536 19708 21548
rect 17819 21508 19708 21536
rect 17819 21505 17831 21508
rect 17773 21499 17831 21505
rect 19702 21496 19708 21508
rect 19760 21496 19766 21548
rect 21818 21536 21824 21548
rect 20088 21508 21824 21536
rect 14461 21471 14519 21477
rect 14461 21437 14473 21471
rect 14507 21437 14519 21471
rect 14461 21431 14519 21437
rect 14553 21471 14611 21477
rect 14553 21437 14565 21471
rect 14599 21437 14611 21471
rect 15010 21468 15016 21480
rect 14971 21440 15016 21468
rect 14553 21431 14611 21437
rect 12268 21372 12322 21400
rect 12366 21372 12572 21400
rect 9858 21332 9864 21344
rect 8260 21304 9864 21332
rect 8260 21292 8266 21304
rect 9858 21292 9864 21304
rect 9916 21292 9922 21344
rect 12294 21332 12322 21372
rect 12434 21332 12440 21344
rect 12294 21304 12440 21332
rect 12434 21292 12440 21304
rect 12492 21292 12498 21344
rect 12544 21332 12572 21372
rect 13998 21360 14004 21412
rect 14056 21400 14062 21412
rect 14568 21400 14596 21431
rect 15010 21428 15016 21440
rect 15068 21428 15074 21480
rect 15473 21471 15531 21477
rect 15473 21437 15485 21471
rect 15519 21437 15531 21471
rect 15473 21431 15531 21437
rect 14056 21372 14596 21400
rect 14056 21360 14062 21372
rect 12802 21332 12808 21344
rect 12544 21304 12808 21332
rect 12802 21292 12808 21304
rect 12860 21332 12866 21344
rect 15488 21332 15516 21431
rect 17678 21428 17684 21480
rect 17736 21468 17742 21480
rect 20088 21477 20116 21508
rect 21818 21496 21824 21508
rect 21876 21496 21882 21548
rect 21910 21496 21916 21548
rect 21968 21536 21974 21548
rect 22557 21539 22615 21545
rect 22557 21536 22569 21539
rect 21968 21508 22569 21536
rect 21968 21496 21974 21508
rect 22557 21505 22569 21508
rect 22603 21505 22615 21539
rect 22557 21499 22615 21505
rect 22646 21496 22652 21548
rect 22704 21536 22710 21548
rect 25608 21536 25636 21644
rect 29454 21632 29460 21644
rect 29512 21632 29518 21684
rect 27246 21564 27252 21616
rect 27304 21604 27310 21616
rect 28445 21607 28503 21613
rect 28445 21604 28457 21607
rect 27304 21576 28457 21604
rect 27304 21564 27310 21576
rect 28445 21573 28457 21576
rect 28491 21573 28503 21607
rect 28445 21567 28503 21573
rect 30561 21607 30619 21613
rect 30561 21573 30573 21607
rect 30607 21573 30619 21607
rect 30561 21567 30619 21573
rect 22704 21508 24624 21536
rect 22704 21496 22710 21508
rect 17957 21471 18015 21477
rect 17957 21468 17969 21471
rect 17736 21440 17969 21468
rect 17736 21428 17742 21440
rect 17957 21437 17969 21440
rect 18003 21437 18015 21471
rect 17957 21431 18015 21437
rect 20073 21471 20131 21477
rect 20073 21437 20085 21471
rect 20119 21437 20131 21471
rect 20073 21431 20131 21437
rect 21453 21471 21511 21477
rect 21453 21437 21465 21471
rect 21499 21437 21511 21471
rect 21453 21431 21511 21437
rect 21637 21471 21695 21477
rect 21637 21437 21649 21471
rect 21683 21468 21695 21471
rect 22922 21468 22928 21480
rect 21683 21440 22928 21468
rect 21683 21437 21695 21440
rect 21637 21431 21695 21437
rect 18690 21360 18696 21412
rect 18748 21400 18754 21412
rect 21468 21400 21496 21431
rect 22922 21428 22928 21440
rect 22980 21428 22986 21480
rect 23017 21471 23075 21477
rect 23017 21437 23029 21471
rect 23063 21468 23075 21471
rect 23566 21468 23572 21480
rect 23063 21440 23572 21468
rect 23063 21437 23075 21440
rect 23017 21431 23075 21437
rect 23566 21428 23572 21440
rect 23624 21428 23630 21480
rect 24596 21477 24624 21508
rect 24688 21508 25636 21536
rect 24581 21471 24639 21477
rect 24581 21437 24593 21471
rect 24627 21437 24639 21471
rect 24581 21431 24639 21437
rect 18748 21372 21496 21400
rect 18748 21360 18754 21372
rect 22462 21360 22468 21412
rect 22520 21400 22526 21412
rect 22695 21403 22753 21409
rect 22695 21400 22707 21403
rect 22520 21372 22707 21400
rect 22520 21360 22526 21372
rect 22695 21369 22707 21372
rect 22741 21369 22753 21403
rect 22695 21363 22753 21369
rect 22833 21403 22891 21409
rect 22833 21369 22845 21403
rect 22879 21400 22891 21403
rect 23106 21400 23112 21412
rect 22879 21372 23112 21400
rect 22879 21369 22891 21372
rect 22833 21363 22891 21369
rect 23106 21360 23112 21372
rect 23164 21400 23170 21412
rect 24688 21400 24716 21508
rect 27062 21496 27068 21548
rect 27120 21536 27126 21548
rect 30576 21536 30604 21567
rect 31202 21536 31208 21548
rect 27120 21508 30420 21536
rect 30576 21508 31208 21536
rect 27120 21496 27126 21508
rect 24854 21468 24860 21480
rect 24815 21440 24860 21468
rect 24854 21428 24860 21440
rect 24912 21428 24918 21480
rect 27982 21468 27988 21480
rect 27943 21440 27988 21468
rect 27982 21428 27988 21440
rect 28040 21428 28046 21480
rect 28166 21428 28172 21480
rect 28224 21468 28230 21480
rect 30392 21477 30420 21508
rect 31202 21496 31208 21508
rect 31260 21536 31266 21548
rect 31386 21536 31392 21548
rect 31260 21508 31392 21536
rect 31260 21496 31266 21508
rect 31386 21496 31392 21508
rect 31444 21536 31450 21548
rect 31481 21539 31539 21545
rect 31481 21536 31493 21539
rect 31444 21508 31493 21536
rect 31444 21496 31450 21508
rect 31481 21505 31493 21508
rect 31527 21505 31539 21539
rect 31481 21499 31539 21505
rect 31665 21539 31723 21545
rect 31665 21505 31677 21539
rect 31711 21536 31723 21539
rect 31846 21536 31852 21548
rect 31711 21508 31852 21536
rect 31711 21505 31723 21508
rect 31665 21499 31723 21505
rect 31846 21496 31852 21508
rect 31904 21536 31910 21548
rect 32950 21536 32956 21548
rect 31904 21508 32956 21536
rect 31904 21496 31910 21508
rect 32950 21496 32956 21508
rect 33008 21496 33014 21548
rect 28261 21471 28319 21477
rect 28261 21468 28273 21471
rect 28224 21440 28273 21468
rect 28224 21428 28230 21440
rect 28261 21437 28273 21440
rect 28307 21437 28319 21471
rect 28261 21431 28319 21437
rect 30377 21471 30435 21477
rect 30377 21437 30389 21471
rect 30423 21437 30435 21471
rect 33594 21468 33600 21480
rect 33555 21440 33600 21468
rect 30377 21431 30435 21437
rect 33594 21428 33600 21440
rect 33652 21428 33658 21480
rect 23164 21372 24716 21400
rect 23164 21360 23170 21372
rect 25314 21360 25320 21412
rect 25372 21400 25378 21412
rect 25685 21403 25743 21409
rect 25685 21400 25697 21403
rect 25372 21372 25697 21400
rect 25372 21360 25378 21372
rect 25685 21369 25697 21372
rect 25731 21369 25743 21403
rect 25685 21363 25743 21369
rect 26418 21360 26424 21412
rect 26476 21400 26482 21412
rect 29181 21403 29239 21409
rect 29181 21400 29193 21403
rect 26476 21372 29193 21400
rect 26476 21360 26482 21372
rect 29181 21369 29193 21372
rect 29227 21369 29239 21403
rect 29181 21363 29239 21369
rect 31757 21403 31815 21409
rect 31757 21369 31769 21403
rect 31803 21400 31815 21403
rect 32214 21400 32220 21412
rect 31803 21372 32220 21400
rect 31803 21369 31815 21372
rect 31757 21363 31815 21369
rect 32214 21360 32220 21372
rect 32272 21360 32278 21412
rect 12860 21304 15516 21332
rect 18141 21335 18199 21341
rect 12860 21292 12866 21304
rect 18141 21301 18153 21335
rect 18187 21332 18199 21335
rect 18506 21332 18512 21344
rect 18187 21304 18512 21332
rect 18187 21301 18199 21304
rect 18141 21295 18199 21301
rect 18506 21292 18512 21304
rect 18564 21292 18570 21344
rect 22922 21292 22928 21344
rect 22980 21332 22986 21344
rect 23934 21332 23940 21344
rect 22980 21304 23940 21332
rect 22980 21292 22986 21304
rect 23934 21292 23940 21304
rect 23992 21332 23998 21344
rect 25480 21335 25538 21341
rect 25480 21332 25492 21335
rect 23992 21304 25492 21332
rect 23992 21292 23998 21304
rect 25480 21301 25492 21304
rect 25526 21332 25538 21335
rect 26142 21332 26148 21344
rect 25526 21304 26148 21332
rect 25526 21301 25538 21304
rect 25480 21295 25538 21301
rect 26142 21292 26148 21304
rect 26200 21292 26206 21344
rect 28994 21292 29000 21344
rect 29052 21332 29058 21344
rect 29089 21335 29147 21341
rect 29089 21332 29101 21335
rect 29052 21304 29101 21332
rect 29052 21292 29058 21304
rect 29089 21301 29101 21304
rect 29135 21301 29147 21335
rect 32122 21332 32128 21344
rect 32083 21304 32128 21332
rect 29089 21295 29147 21301
rect 32122 21292 32128 21304
rect 32180 21292 32186 21344
rect 33410 21332 33416 21344
rect 33371 21304 33416 21332
rect 33410 21292 33416 21304
rect 33468 21292 33474 21344
rect 1104 21242 34316 21264
rect 1104 21190 12052 21242
rect 12104 21190 12116 21242
rect 12168 21190 12180 21242
rect 12232 21190 12244 21242
rect 12296 21190 23123 21242
rect 23175 21190 23187 21242
rect 23239 21190 23251 21242
rect 23303 21190 23315 21242
rect 23367 21190 34316 21242
rect 1104 21168 34316 21190
rect 4338 21088 4344 21140
rect 4396 21128 4402 21140
rect 4985 21131 5043 21137
rect 4985 21128 4997 21131
rect 4396 21100 4997 21128
rect 4396 21088 4402 21100
rect 4985 21097 4997 21100
rect 5031 21097 5043 21131
rect 6914 21128 6920 21140
rect 4985 21091 5043 21097
rect 5184 21100 6920 21128
rect 2961 21063 3019 21069
rect 2961 21029 2973 21063
rect 3007 21060 3019 21063
rect 3970 21060 3976 21072
rect 3007 21032 3976 21060
rect 3007 21029 3019 21032
rect 2961 21023 3019 21029
rect 3970 21020 3976 21032
rect 4028 21020 4034 21072
rect 3142 20992 3148 21004
rect 3103 20964 3148 20992
rect 3142 20952 3148 20964
rect 3200 20952 3206 21004
rect 3237 20995 3295 21001
rect 3237 20961 3249 20995
rect 3283 20961 3295 20995
rect 3237 20955 3295 20961
rect 3252 20924 3280 20955
rect 3326 20952 3332 21004
rect 3384 20992 3390 21004
rect 5184 21001 5212 21100
rect 6914 21088 6920 21100
rect 6972 21088 6978 21140
rect 7282 21128 7288 21140
rect 7243 21100 7288 21128
rect 7282 21088 7288 21100
rect 7340 21088 7346 21140
rect 8662 21088 8668 21140
rect 8720 21128 8726 21140
rect 11422 21128 11428 21140
rect 8720 21100 10364 21128
rect 11383 21100 11428 21128
rect 8720 21088 8726 21100
rect 6457 21063 6515 21069
rect 6457 21060 6469 21063
rect 5736 21032 6469 21060
rect 4249 20995 4307 21001
rect 4249 20992 4261 20995
rect 3384 20964 4261 20992
rect 3384 20952 3390 20964
rect 4249 20961 4261 20964
rect 4295 20961 4307 20995
rect 4249 20955 4307 20961
rect 5169 20995 5227 21001
rect 5169 20961 5181 20995
rect 5215 20961 5227 20995
rect 5169 20955 5227 20961
rect 5353 20995 5411 21001
rect 5353 20961 5365 20995
rect 5399 20992 5411 20995
rect 5442 20992 5448 21004
rect 5399 20964 5448 20992
rect 5399 20961 5411 20964
rect 5353 20955 5411 20961
rect 5442 20952 5448 20964
rect 5500 20952 5506 21004
rect 5534 20952 5540 21004
rect 5592 20992 5598 21004
rect 5736 21001 5764 21032
rect 6457 21029 6469 21032
rect 6503 21029 6515 21063
rect 8202 21060 8208 21072
rect 8163 21032 8208 21060
rect 6457 21023 6515 21029
rect 8202 21020 8208 21032
rect 8260 21020 8266 21072
rect 8297 21063 8355 21069
rect 8297 21029 8309 21063
rect 8343 21060 8355 21063
rect 9306 21060 9312 21072
rect 8343 21032 9312 21060
rect 8343 21029 8355 21032
rect 8297 21023 8355 21029
rect 9306 21020 9312 21032
rect 9364 21020 9370 21072
rect 9493 21063 9551 21069
rect 9493 21029 9505 21063
rect 9539 21060 9551 21063
rect 9582 21060 9588 21072
rect 9539 21032 9588 21060
rect 9539 21029 9551 21032
rect 9493 21023 9551 21029
rect 9582 21020 9588 21032
rect 9640 21020 9646 21072
rect 9677 21063 9735 21069
rect 9677 21029 9689 21063
rect 9723 21060 9735 21063
rect 9858 21060 9864 21072
rect 9723 21032 9864 21060
rect 9723 21029 9735 21032
rect 9677 21023 9735 21029
rect 9858 21020 9864 21032
rect 9916 21020 9922 21072
rect 5721 20995 5779 21001
rect 5721 20992 5733 20995
rect 5592 20964 5733 20992
rect 5592 20952 5598 20964
rect 5721 20961 5733 20964
rect 5767 20961 5779 20995
rect 6362 20992 6368 21004
rect 6323 20964 6368 20992
rect 5721 20955 5779 20961
rect 6362 20952 6368 20964
rect 6420 20952 6426 21004
rect 7006 20952 7012 21004
rect 7064 20992 7070 21004
rect 10336 21001 10364 21100
rect 11422 21088 11428 21100
rect 11480 21088 11486 21140
rect 11882 21088 11888 21140
rect 11940 21128 11946 21140
rect 11940 21100 12020 21128
rect 11940 21088 11946 21100
rect 11992 21069 12020 21100
rect 15010 21088 15016 21140
rect 15068 21128 15074 21140
rect 15841 21131 15899 21137
rect 15841 21128 15853 21131
rect 15068 21100 15853 21128
rect 15068 21088 15074 21100
rect 15841 21097 15853 21100
rect 15887 21097 15899 21131
rect 15841 21091 15899 21097
rect 17402 21088 17408 21140
rect 17460 21128 17466 21140
rect 17678 21128 17684 21140
rect 17460 21100 17684 21128
rect 17460 21088 17466 21100
rect 17678 21088 17684 21100
rect 17736 21088 17742 21140
rect 33410 21128 33416 21140
rect 22066 21100 33416 21128
rect 11977 21063 12035 21069
rect 11977 21029 11989 21063
rect 12023 21029 12035 21063
rect 12802 21060 12808 21072
rect 11977 21023 12035 21029
rect 12360 21032 12808 21060
rect 7193 20995 7251 21001
rect 7193 20992 7205 20995
rect 7064 20964 7205 20992
rect 7064 20952 7070 20964
rect 7193 20961 7205 20964
rect 7239 20961 7251 20995
rect 7193 20955 7251 20961
rect 8113 20995 8171 21001
rect 8113 20961 8125 20995
rect 8159 20961 8171 20995
rect 8113 20955 8171 20961
rect 8435 20995 8493 21001
rect 8435 20961 8447 20995
rect 8481 20992 8493 20995
rect 10321 20995 10379 21001
rect 8481 20964 9628 20992
rect 8481 20961 8493 20964
rect 8435 20955 8493 20961
rect 4430 20924 4436 20936
rect 3252 20896 4436 20924
rect 4430 20884 4436 20896
rect 4488 20884 4494 20936
rect 4522 20884 4528 20936
rect 4580 20924 4586 20936
rect 4893 20927 4951 20933
rect 4893 20924 4905 20927
rect 4580 20896 4905 20924
rect 4580 20884 4586 20896
rect 4893 20893 4905 20896
rect 4939 20893 4951 20927
rect 4893 20887 4951 20893
rect 5629 20927 5687 20933
rect 5629 20893 5641 20927
rect 5675 20893 5687 20927
rect 5629 20887 5687 20893
rect 2958 20856 2964 20868
rect 2919 20828 2964 20856
rect 2958 20816 2964 20828
rect 3016 20816 3022 20868
rect 4341 20859 4399 20865
rect 4341 20825 4353 20859
rect 4387 20856 4399 20859
rect 4614 20856 4620 20868
rect 4387 20828 4620 20856
rect 4387 20825 4399 20828
rect 4341 20819 4399 20825
rect 4614 20816 4620 20828
rect 4672 20856 4678 20868
rect 5644 20856 5672 20887
rect 4672 20828 5672 20856
rect 8128 20856 8156 20955
rect 9600 20936 9628 20964
rect 10321 20961 10333 20995
rect 10367 20961 10379 20995
rect 10321 20955 10379 20961
rect 10505 20995 10563 21001
rect 10505 20961 10517 20995
rect 10551 20992 10563 20995
rect 10962 20992 10968 21004
rect 10551 20964 10968 20992
rect 10551 20961 10563 20964
rect 10505 20955 10563 20961
rect 8202 20884 8208 20936
rect 8260 20924 8266 20936
rect 8573 20927 8631 20933
rect 8573 20924 8585 20927
rect 8260 20896 8585 20924
rect 8260 20884 8266 20896
rect 8573 20893 8585 20896
rect 8619 20893 8631 20927
rect 8573 20887 8631 20893
rect 9582 20884 9588 20936
rect 9640 20884 9646 20936
rect 9766 20884 9772 20936
rect 9824 20924 9830 20936
rect 10520 20924 10548 20955
rect 10962 20952 10968 20964
rect 11020 20952 11026 21004
rect 11241 20995 11299 21001
rect 11241 20961 11253 20995
rect 11287 20961 11299 20995
rect 11241 20955 11299 20961
rect 11425 20995 11483 21001
rect 11425 20961 11437 20995
rect 11471 20961 11483 20995
rect 11882 20992 11888 21004
rect 11843 20964 11888 20992
rect 11425 20955 11483 20961
rect 9824 20896 10548 20924
rect 9824 20884 9830 20896
rect 10321 20859 10379 20865
rect 10321 20856 10333 20859
rect 8128 20828 10333 20856
rect 4672 20816 4678 20828
rect 10321 20825 10333 20828
rect 10367 20825 10379 20859
rect 10321 20819 10379 20825
rect 3970 20748 3976 20800
rect 4028 20788 4034 20800
rect 6362 20788 6368 20800
rect 4028 20760 6368 20788
rect 4028 20748 4034 20760
rect 6362 20748 6368 20760
rect 6420 20748 6426 20800
rect 7929 20791 7987 20797
rect 7929 20757 7941 20791
rect 7975 20788 7987 20791
rect 8386 20788 8392 20800
rect 7975 20760 8392 20788
rect 7975 20757 7987 20760
rect 7929 20751 7987 20757
rect 8386 20748 8392 20760
rect 8444 20748 8450 20800
rect 9861 20791 9919 20797
rect 9861 20757 9873 20791
rect 9907 20788 9919 20791
rect 10502 20788 10508 20800
rect 9907 20760 10508 20788
rect 9907 20757 9919 20760
rect 9861 20751 9919 20757
rect 10502 20748 10508 20760
rect 10560 20748 10566 20800
rect 11256 20788 11284 20955
rect 11440 20924 11468 20955
rect 11882 20952 11888 20964
rect 11940 20952 11946 21004
rect 12360 21001 12388 21032
rect 12802 21020 12808 21032
rect 12860 21020 12866 21072
rect 22066 21060 22094 21100
rect 33410 21088 33416 21100
rect 33468 21088 33474 21140
rect 22462 21060 22468 21072
rect 15580 21032 22094 21060
rect 22423 21032 22468 21060
rect 12345 20995 12403 21001
rect 12345 20961 12357 20995
rect 12391 20961 12403 20995
rect 12345 20955 12403 20961
rect 12526 20952 12532 21004
rect 12584 20992 12590 21004
rect 12713 20995 12771 21001
rect 12713 20992 12725 20995
rect 12584 20964 12725 20992
rect 12584 20952 12590 20964
rect 12713 20961 12725 20964
rect 12759 20961 12771 20995
rect 12713 20955 12771 20961
rect 14550 20952 14556 21004
rect 14608 20992 14614 21004
rect 15013 20995 15071 21001
rect 15013 20992 15025 20995
rect 14608 20964 15025 20992
rect 14608 20952 14614 20964
rect 15013 20961 15025 20964
rect 15059 20961 15071 20995
rect 15013 20955 15071 20961
rect 15102 20952 15108 21004
rect 15160 20992 15166 21004
rect 15580 20992 15608 21032
rect 22462 21020 22468 21032
rect 22520 21020 22526 21072
rect 24026 21060 24032 21072
rect 23987 21032 24032 21060
rect 24026 21020 24032 21032
rect 24084 21020 24090 21072
rect 24854 21020 24860 21072
rect 24912 21060 24918 21072
rect 25777 21063 25835 21069
rect 25777 21060 25789 21063
rect 24912 21032 25789 21060
rect 24912 21020 24918 21032
rect 25777 21029 25789 21032
rect 25823 21060 25835 21063
rect 27430 21060 27436 21072
rect 25823 21032 27436 21060
rect 25823 21029 25835 21032
rect 25777 21023 25835 21029
rect 27430 21020 27436 21032
rect 27488 21020 27494 21072
rect 32122 21060 32128 21072
rect 32083 21032 32128 21060
rect 32122 21020 32128 21032
rect 32180 21020 32186 21072
rect 32582 21020 32588 21072
rect 32640 21020 32646 21072
rect 16574 21001 16580 21004
rect 15160 20964 15608 20992
rect 15160 20952 15166 20964
rect 16568 20955 16580 21001
rect 16632 20992 16638 21004
rect 18690 20992 18696 21004
rect 16632 20964 16668 20992
rect 18651 20964 18696 20992
rect 16574 20952 16580 20955
rect 16632 20952 16638 20964
rect 18690 20952 18696 20964
rect 18748 20952 18754 21004
rect 20346 20992 20352 21004
rect 20307 20964 20352 20992
rect 20346 20952 20352 20964
rect 20404 20952 20410 21004
rect 22370 20992 22376 21004
rect 22331 20964 22376 20992
rect 22370 20952 22376 20964
rect 22428 20952 22434 21004
rect 22557 20995 22615 21001
rect 22557 20961 22569 20995
rect 22603 20992 22615 20995
rect 22738 20992 22744 21004
rect 22603 20964 22744 20992
rect 22603 20961 22615 20964
rect 22557 20955 22615 20961
rect 22738 20952 22744 20964
rect 22796 20952 22802 21004
rect 23293 20995 23351 21001
rect 23293 20961 23305 20995
rect 23339 20961 23351 20995
rect 23293 20955 23351 20961
rect 23477 20995 23535 21001
rect 23477 20961 23489 20995
rect 23523 20961 23535 20995
rect 23477 20955 23535 20961
rect 12250 20924 12256 20936
rect 11440 20896 12256 20924
rect 12250 20884 12256 20896
rect 12308 20884 12314 20936
rect 12434 20924 12440 20936
rect 12395 20896 12440 20924
rect 12434 20884 12440 20896
rect 12492 20884 12498 20936
rect 12621 20927 12679 20933
rect 12621 20893 12633 20927
rect 12667 20893 12679 20927
rect 14918 20924 14924 20936
rect 14879 20896 14924 20924
rect 12621 20887 12679 20893
rect 12636 20788 12664 20887
rect 14918 20884 14924 20896
rect 14976 20884 14982 20936
rect 16298 20924 16304 20936
rect 16259 20896 16304 20924
rect 16298 20884 16304 20896
rect 16356 20884 16362 20936
rect 18969 20927 19027 20933
rect 18969 20893 18981 20927
rect 19015 20924 19027 20927
rect 19426 20924 19432 20936
rect 19015 20896 19432 20924
rect 19015 20893 19027 20896
rect 18969 20887 19027 20893
rect 19426 20884 19432 20896
rect 19484 20884 19490 20936
rect 20257 20927 20315 20933
rect 20257 20893 20269 20927
rect 20303 20924 20315 20927
rect 20990 20924 20996 20936
rect 20303 20896 20996 20924
rect 20303 20893 20315 20896
rect 20257 20887 20315 20893
rect 20990 20884 20996 20896
rect 21048 20884 21054 20936
rect 22388 20924 22416 20952
rect 23308 20924 23336 20955
rect 22388 20896 23336 20924
rect 23492 20924 23520 20955
rect 23750 20952 23756 21004
rect 23808 20992 23814 21004
rect 23934 20992 23940 21004
rect 23808 20964 23940 20992
rect 23808 20952 23814 20964
rect 23934 20952 23940 20964
rect 23992 20952 23998 21004
rect 25498 20952 25504 21004
rect 25556 20992 25562 21004
rect 25593 20995 25651 21001
rect 25593 20992 25605 20995
rect 25556 20964 25605 20992
rect 25556 20952 25562 20964
rect 25593 20961 25605 20964
rect 25639 20992 25651 20995
rect 26142 20992 26148 21004
rect 25639 20964 26148 20992
rect 25639 20961 25651 20964
rect 25593 20955 25651 20961
rect 26142 20952 26148 20964
rect 26200 20952 26206 21004
rect 26510 20992 26516 21004
rect 26471 20964 26516 20992
rect 26510 20952 26516 20964
rect 26568 20952 26574 21004
rect 27246 20992 27252 21004
rect 27207 20964 27252 20992
rect 27246 20952 27252 20964
rect 27304 20952 27310 21004
rect 29086 20992 29092 21004
rect 29144 21001 29150 21004
rect 29056 20964 29092 20992
rect 29086 20952 29092 20964
rect 29144 20955 29156 21001
rect 30834 20992 30840 21004
rect 30795 20964 30840 20992
rect 29144 20952 29150 20955
rect 30834 20952 30840 20964
rect 30892 20952 30898 21004
rect 25222 20924 25228 20936
rect 23492 20896 25228 20924
rect 25222 20884 25228 20896
rect 25280 20884 25286 20936
rect 25314 20884 25320 20936
rect 25372 20924 25378 20936
rect 25409 20927 25467 20933
rect 25409 20924 25421 20927
rect 25372 20896 25421 20924
rect 25372 20884 25378 20896
rect 25409 20893 25421 20896
rect 25455 20893 25467 20927
rect 25409 20887 25467 20893
rect 26418 20884 26424 20936
rect 26476 20924 26482 20936
rect 26476 20896 27108 20924
rect 26476 20884 26482 20896
rect 18877 20859 18935 20865
rect 18877 20825 18889 20859
rect 18923 20856 18935 20859
rect 19058 20856 19064 20868
rect 18923 20828 19064 20856
rect 18923 20825 18935 20828
rect 18877 20819 18935 20825
rect 19058 20816 19064 20828
rect 19116 20816 19122 20868
rect 27080 20865 27108 20896
rect 29362 20884 29368 20936
rect 29420 20924 29426 20936
rect 29822 20924 29828 20936
rect 29420 20896 29828 20924
rect 29420 20884 29426 20896
rect 29822 20884 29828 20896
rect 29880 20884 29886 20936
rect 30929 20927 30987 20933
rect 30929 20893 30941 20927
rect 30975 20893 30987 20927
rect 30929 20887 30987 20893
rect 31113 20927 31171 20933
rect 31113 20893 31125 20927
rect 31159 20924 31171 20927
rect 31202 20924 31208 20936
rect 31159 20896 31208 20924
rect 31159 20893 31171 20896
rect 31113 20887 31171 20893
rect 27065 20859 27123 20865
rect 27065 20825 27077 20859
rect 27111 20825 27123 20859
rect 30944 20856 30972 20887
rect 31202 20884 31208 20896
rect 31260 20884 31266 20936
rect 31754 20884 31760 20936
rect 31812 20924 31818 20936
rect 31849 20927 31907 20933
rect 31849 20924 31861 20927
rect 31812 20896 31861 20924
rect 31812 20884 31818 20896
rect 31849 20893 31861 20896
rect 31895 20893 31907 20927
rect 32214 20924 32220 20936
rect 31849 20887 31907 20893
rect 31956 20896 32220 20924
rect 31956 20856 31984 20896
rect 32214 20884 32220 20896
rect 32272 20924 32278 20936
rect 33597 20927 33655 20933
rect 33597 20924 33609 20927
rect 32272 20896 33609 20924
rect 32272 20884 32278 20896
rect 33597 20893 33609 20896
rect 33643 20893 33655 20927
rect 33597 20887 33655 20893
rect 30944 20828 31984 20856
rect 27065 20819 27123 20825
rect 12894 20788 12900 20800
rect 11256 20760 12900 20788
rect 12894 20748 12900 20760
rect 12952 20748 12958 20800
rect 18322 20748 18328 20800
rect 18380 20788 18386 20800
rect 18509 20791 18567 20797
rect 18509 20788 18521 20791
rect 18380 20760 18521 20788
rect 18380 20748 18386 20760
rect 18509 20757 18521 20760
rect 18555 20757 18567 20791
rect 18509 20751 18567 20757
rect 18966 20748 18972 20800
rect 19024 20788 19030 20800
rect 19981 20791 20039 20797
rect 19981 20788 19993 20791
rect 19024 20760 19993 20788
rect 19024 20748 19030 20760
rect 19981 20757 19993 20760
rect 20027 20757 20039 20791
rect 20162 20788 20168 20800
rect 20123 20760 20168 20788
rect 19981 20751 20039 20757
rect 20162 20748 20168 20760
rect 20220 20748 20226 20800
rect 23293 20791 23351 20797
rect 23293 20757 23305 20791
rect 23339 20788 23351 20791
rect 23934 20788 23940 20800
rect 23339 20760 23940 20788
rect 23339 20757 23351 20760
rect 23293 20751 23351 20757
rect 23934 20748 23940 20760
rect 23992 20748 23998 20800
rect 26421 20791 26479 20797
rect 26421 20757 26433 20791
rect 26467 20788 26479 20791
rect 26602 20788 26608 20800
rect 26467 20760 26608 20788
rect 26467 20757 26479 20760
rect 26421 20751 26479 20757
rect 26602 20748 26608 20760
rect 26660 20748 26666 20800
rect 27614 20748 27620 20800
rect 27672 20788 27678 20800
rect 27985 20791 28043 20797
rect 27985 20788 27997 20791
rect 27672 20760 27997 20788
rect 27672 20748 27678 20760
rect 27985 20757 27997 20760
rect 28031 20757 28043 20791
rect 30466 20788 30472 20800
rect 30427 20760 30472 20788
rect 27985 20751 28043 20757
rect 30466 20748 30472 20760
rect 30524 20748 30530 20800
rect 1104 20698 34316 20720
rect 1104 20646 6517 20698
rect 6569 20646 6581 20698
rect 6633 20646 6645 20698
rect 6697 20646 6709 20698
rect 6761 20646 17588 20698
rect 17640 20646 17652 20698
rect 17704 20646 17716 20698
rect 17768 20646 17780 20698
rect 17832 20646 28658 20698
rect 28710 20646 28722 20698
rect 28774 20646 28786 20698
rect 28838 20646 28850 20698
rect 28902 20646 34316 20698
rect 1104 20624 34316 20646
rect 2961 20587 3019 20593
rect 2961 20553 2973 20587
rect 3007 20584 3019 20587
rect 3142 20584 3148 20596
rect 3007 20556 3148 20584
rect 3007 20553 3019 20556
rect 2961 20547 3019 20553
rect 3142 20544 3148 20556
rect 3200 20544 3206 20596
rect 3326 20584 3332 20596
rect 3287 20556 3332 20584
rect 3326 20544 3332 20556
rect 3384 20544 3390 20596
rect 3973 20587 4031 20593
rect 3973 20553 3985 20587
rect 4019 20584 4031 20587
rect 4062 20584 4068 20596
rect 4019 20556 4068 20584
rect 4019 20553 4031 20556
rect 3973 20547 4031 20553
rect 4062 20544 4068 20556
rect 4120 20544 4126 20596
rect 6914 20584 6920 20596
rect 6875 20556 6920 20584
rect 6914 20544 6920 20556
rect 6972 20584 6978 20596
rect 8202 20584 8208 20596
rect 6972 20556 8208 20584
rect 6972 20544 6978 20556
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 9674 20544 9680 20596
rect 9732 20584 9738 20596
rect 10505 20587 10563 20593
rect 10505 20584 10517 20587
rect 9732 20556 10517 20584
rect 9732 20544 9738 20556
rect 10505 20553 10517 20556
rect 10551 20553 10563 20587
rect 10505 20547 10563 20553
rect 10965 20587 11023 20593
rect 10965 20553 10977 20587
rect 11011 20584 11023 20587
rect 11882 20584 11888 20596
rect 11011 20556 11888 20584
rect 11011 20553 11023 20556
rect 10965 20547 11023 20553
rect 11882 20544 11888 20556
rect 11940 20544 11946 20596
rect 12253 20587 12311 20593
rect 12253 20553 12265 20587
rect 12299 20584 12311 20587
rect 12342 20584 12348 20596
rect 12299 20556 12348 20584
rect 12299 20553 12311 20556
rect 12253 20547 12311 20553
rect 12342 20544 12348 20556
rect 12400 20544 12406 20596
rect 19426 20584 19432 20596
rect 19339 20556 19432 20584
rect 19426 20544 19432 20556
rect 19484 20584 19490 20596
rect 20162 20584 20168 20596
rect 19484 20556 20168 20584
rect 19484 20544 19490 20556
rect 20162 20544 20168 20556
rect 20220 20544 20226 20596
rect 23842 20544 23848 20596
rect 23900 20584 23906 20596
rect 24762 20584 24768 20596
rect 23900 20556 24768 20584
rect 23900 20544 23906 20556
rect 24762 20544 24768 20556
rect 24820 20544 24826 20596
rect 25958 20584 25964 20596
rect 25919 20556 25964 20584
rect 25958 20544 25964 20556
rect 26016 20544 26022 20596
rect 26050 20544 26056 20596
rect 26108 20584 26114 20596
rect 26605 20587 26663 20593
rect 26605 20584 26617 20587
rect 26108 20556 26617 20584
rect 26108 20544 26114 20556
rect 26605 20553 26617 20556
rect 26651 20553 26663 20587
rect 26605 20547 26663 20553
rect 28077 20587 28135 20593
rect 28077 20553 28089 20587
rect 28123 20584 28135 20587
rect 29086 20584 29092 20596
rect 28123 20556 29092 20584
rect 28123 20553 28135 20556
rect 28077 20547 28135 20553
rect 29086 20544 29092 20556
rect 29144 20544 29150 20596
rect 30834 20544 30840 20596
rect 30892 20584 30898 20596
rect 31297 20587 31355 20593
rect 31297 20584 31309 20587
rect 30892 20556 31309 20584
rect 30892 20544 30898 20556
rect 31297 20553 31309 20556
rect 31343 20553 31355 20587
rect 31297 20547 31355 20553
rect 13446 20516 13452 20528
rect 10704 20488 13452 20516
rect 1762 20448 1768 20460
rect 1723 20420 1768 20448
rect 1762 20408 1768 20420
rect 1820 20408 1826 20460
rect 3421 20451 3479 20457
rect 3421 20417 3433 20451
rect 3467 20448 3479 20451
rect 3970 20448 3976 20460
rect 3467 20420 3976 20448
rect 3467 20417 3479 20420
rect 3421 20411 3479 20417
rect 3970 20408 3976 20420
rect 4028 20408 4034 20460
rect 8386 20448 8392 20460
rect 8347 20420 8392 20448
rect 8386 20408 8392 20420
rect 8444 20408 8450 20460
rect 8665 20451 8723 20457
rect 8665 20417 8677 20451
rect 8711 20448 8723 20451
rect 9398 20448 9404 20460
rect 8711 20420 9404 20448
rect 8711 20417 8723 20420
rect 8665 20411 8723 20417
rect 9398 20408 9404 20420
rect 9456 20408 9462 20460
rect 3145 20383 3203 20389
rect 3145 20349 3157 20383
rect 3191 20349 3203 20383
rect 3878 20380 3884 20392
rect 3839 20352 3884 20380
rect 3145 20343 3203 20349
rect 1946 20312 1952 20324
rect 1907 20284 1952 20312
rect 1946 20272 1952 20284
rect 2004 20272 2010 20324
rect 3160 20312 3188 20343
rect 3878 20340 3884 20352
rect 3936 20340 3942 20392
rect 4798 20340 4804 20392
rect 4856 20380 4862 20392
rect 5077 20383 5135 20389
rect 5077 20380 5089 20383
rect 4856 20352 5089 20380
rect 4856 20340 4862 20352
rect 5077 20349 5089 20352
rect 5123 20349 5135 20383
rect 5077 20343 5135 20349
rect 5442 20340 5448 20392
rect 5500 20380 5506 20392
rect 5537 20383 5595 20389
rect 5537 20380 5549 20383
rect 5500 20352 5549 20380
rect 5500 20340 5506 20352
rect 5537 20349 5549 20352
rect 5583 20349 5595 20383
rect 5718 20380 5724 20392
rect 5679 20352 5724 20380
rect 5537 20343 5595 20349
rect 5718 20340 5724 20352
rect 5776 20340 5782 20392
rect 9585 20383 9643 20389
rect 9585 20349 9597 20383
rect 9631 20380 9643 20383
rect 9950 20380 9956 20392
rect 9631 20352 9956 20380
rect 9631 20349 9643 20352
rect 9585 20343 9643 20349
rect 9950 20340 9956 20352
rect 10008 20380 10014 20392
rect 10502 20380 10508 20392
rect 10008 20352 10364 20380
rect 10463 20352 10508 20380
rect 10008 20340 10014 20352
rect 5629 20315 5687 20321
rect 5629 20312 5641 20315
rect 3160 20284 5641 20312
rect 5629 20281 5641 20284
rect 5675 20281 5687 20315
rect 5629 20275 5687 20281
rect 7006 20272 7012 20324
rect 7064 20312 7070 20324
rect 7064 20284 7222 20312
rect 7064 20272 7070 20284
rect 8938 20272 8944 20324
rect 8996 20312 9002 20324
rect 9677 20315 9735 20321
rect 9677 20312 9689 20315
rect 8996 20284 9689 20312
rect 8996 20272 9002 20284
rect 9677 20281 9689 20284
rect 9723 20281 9735 20315
rect 9677 20275 9735 20281
rect 4985 20247 5043 20253
rect 4985 20213 4997 20247
rect 5031 20244 5043 20247
rect 5074 20244 5080 20256
rect 5031 20216 5080 20244
rect 5031 20213 5043 20216
rect 4985 20207 5043 20213
rect 5074 20204 5080 20216
rect 5132 20204 5138 20256
rect 10336 20244 10364 20352
rect 10502 20340 10508 20352
rect 10560 20340 10566 20392
rect 10704 20389 10732 20488
rect 13446 20476 13452 20488
rect 13504 20476 13510 20528
rect 13538 20476 13544 20528
rect 13596 20516 13602 20528
rect 17405 20519 17463 20525
rect 17405 20516 17417 20519
rect 13596 20488 17417 20516
rect 13596 20476 13602 20488
rect 17405 20485 17417 20488
rect 17451 20485 17463 20519
rect 27246 20516 27252 20528
rect 17405 20479 17463 20485
rect 22066 20488 27252 20516
rect 12176 20420 16068 20448
rect 10689 20383 10747 20389
rect 10689 20349 10701 20383
rect 10735 20349 10747 20383
rect 10689 20343 10747 20349
rect 10781 20383 10839 20389
rect 10781 20349 10793 20383
rect 10827 20349 10839 20383
rect 11054 20380 11060 20392
rect 11015 20352 11060 20380
rect 10781 20343 10839 20349
rect 10796 20312 10824 20343
rect 11054 20340 11060 20352
rect 11112 20340 11118 20392
rect 11330 20340 11336 20392
rect 11388 20380 11394 20392
rect 12176 20389 12204 20420
rect 12161 20383 12219 20389
rect 12161 20380 12173 20383
rect 11388 20352 12173 20380
rect 11388 20340 11394 20352
rect 12161 20349 12173 20352
rect 12207 20349 12219 20383
rect 12161 20343 12219 20349
rect 12345 20383 12403 20389
rect 12345 20349 12357 20383
rect 12391 20380 12403 20383
rect 12526 20380 12532 20392
rect 12391 20352 12532 20380
rect 12391 20349 12403 20352
rect 12345 20343 12403 20349
rect 12526 20340 12532 20352
rect 12584 20340 12590 20392
rect 13170 20340 13176 20392
rect 13228 20380 13234 20392
rect 13357 20383 13415 20389
rect 13357 20380 13369 20383
rect 13228 20352 13369 20380
rect 13228 20340 13234 20352
rect 13357 20349 13369 20352
rect 13403 20349 13415 20383
rect 13357 20343 13415 20349
rect 13541 20383 13599 20389
rect 13541 20349 13553 20383
rect 13587 20380 13599 20383
rect 13630 20380 13636 20392
rect 13587 20352 13636 20380
rect 13587 20349 13599 20352
rect 13541 20343 13599 20349
rect 13630 20340 13636 20352
rect 13688 20340 13694 20392
rect 13998 20380 14004 20392
rect 13959 20352 14004 20380
rect 13998 20340 14004 20352
rect 14056 20340 14062 20392
rect 14185 20383 14243 20389
rect 14185 20349 14197 20383
rect 14231 20349 14243 20383
rect 14185 20343 14243 20349
rect 10962 20312 10968 20324
rect 10796 20284 10968 20312
rect 10962 20272 10968 20284
rect 11020 20272 11026 20324
rect 12434 20272 12440 20324
rect 12492 20312 12498 20324
rect 13262 20312 13268 20324
rect 12492 20284 13268 20312
rect 12492 20272 12498 20284
rect 13262 20272 13268 20284
rect 13320 20312 13326 20324
rect 14200 20312 14228 20343
rect 15838 20312 15844 20324
rect 13320 20284 14228 20312
rect 15799 20284 15844 20312
rect 13320 20272 13326 20284
rect 15838 20272 15844 20284
rect 15896 20272 15902 20324
rect 16040 20321 16068 20420
rect 16298 20408 16304 20460
rect 16356 20448 16362 20460
rect 18049 20451 18107 20457
rect 18049 20448 18061 20451
rect 16356 20420 18061 20448
rect 16356 20408 16362 20420
rect 18049 20417 18061 20420
rect 18095 20417 18107 20451
rect 18049 20411 18107 20417
rect 17310 20380 17316 20392
rect 17271 20352 17316 20380
rect 17310 20340 17316 20352
rect 17368 20340 17374 20392
rect 17402 20340 17408 20392
rect 17460 20380 17466 20392
rect 18322 20389 18328 20392
rect 17497 20383 17555 20389
rect 17497 20380 17509 20383
rect 17460 20352 17509 20380
rect 17460 20340 17466 20352
rect 17497 20349 17509 20352
rect 17543 20349 17555 20383
rect 18316 20380 18328 20389
rect 18283 20352 18328 20380
rect 17497 20343 17555 20349
rect 18316 20343 18328 20352
rect 18322 20340 18328 20343
rect 18380 20340 18386 20392
rect 20717 20383 20775 20389
rect 20717 20349 20729 20383
rect 20763 20380 20775 20383
rect 20990 20380 20996 20392
rect 20763 20352 20996 20380
rect 20763 20349 20775 20352
rect 20717 20343 20775 20349
rect 20990 20340 20996 20352
rect 21048 20340 21054 20392
rect 21269 20383 21327 20389
rect 21269 20349 21281 20383
rect 21315 20380 21327 20383
rect 22066 20380 22094 20488
rect 27246 20476 27252 20488
rect 27304 20476 27310 20528
rect 22186 20408 22192 20460
rect 22244 20448 22250 20460
rect 22554 20448 22560 20460
rect 22244 20420 22560 20448
rect 22244 20408 22250 20420
rect 22554 20408 22560 20420
rect 22612 20448 22618 20460
rect 22612 20420 23888 20448
rect 22612 20408 22618 20420
rect 23014 20380 23020 20392
rect 21315 20352 22094 20380
rect 22975 20352 23020 20380
rect 21315 20349 21327 20352
rect 21269 20343 21327 20349
rect 23014 20340 23020 20352
rect 23072 20340 23078 20392
rect 23474 20380 23480 20392
rect 23435 20352 23480 20380
rect 23474 20340 23480 20352
rect 23532 20340 23538 20392
rect 23750 20380 23756 20392
rect 23711 20352 23756 20380
rect 23750 20340 23756 20352
rect 23808 20340 23814 20392
rect 23860 20380 23888 20420
rect 23934 20408 23940 20460
rect 23992 20448 23998 20460
rect 23992 20420 25176 20448
rect 23992 20408 23998 20420
rect 25148 20389 25176 20420
rect 28258 20408 28264 20460
rect 28316 20448 28322 20460
rect 28629 20451 28687 20457
rect 28629 20448 28641 20451
rect 28316 20420 28641 20448
rect 28316 20408 28322 20420
rect 28629 20417 28641 20420
rect 28675 20448 28687 20451
rect 28994 20448 29000 20460
rect 28675 20420 29000 20448
rect 28675 20417 28687 20420
rect 28629 20411 28687 20417
rect 28994 20408 29000 20420
rect 29052 20408 29058 20460
rect 29825 20451 29883 20457
rect 29825 20417 29837 20451
rect 29871 20448 29883 20451
rect 30466 20448 30472 20460
rect 29871 20420 30472 20448
rect 29871 20417 29883 20420
rect 29825 20411 29883 20417
rect 30466 20408 30472 20420
rect 30524 20408 30530 20460
rect 24673 20383 24731 20389
rect 24673 20380 24685 20383
rect 23860 20352 24685 20380
rect 24673 20349 24685 20352
rect 24719 20349 24731 20383
rect 24673 20343 24731 20349
rect 25041 20383 25099 20389
rect 25041 20349 25053 20383
rect 25087 20349 25099 20383
rect 25041 20343 25099 20349
rect 25133 20383 25191 20389
rect 25133 20349 25145 20383
rect 25179 20349 25191 20383
rect 25133 20343 25191 20349
rect 16025 20315 16083 20321
rect 16025 20281 16037 20315
rect 16071 20312 16083 20315
rect 16114 20312 16120 20324
rect 16071 20284 16120 20312
rect 16071 20281 16083 20284
rect 16025 20275 16083 20281
rect 16114 20272 16120 20284
rect 16172 20272 16178 20324
rect 16758 20272 16764 20324
rect 16816 20312 16822 20324
rect 17420 20312 17448 20340
rect 22830 20312 22836 20324
rect 16816 20284 17448 20312
rect 22791 20284 22836 20312
rect 16816 20272 16822 20284
rect 22830 20272 22836 20284
rect 22888 20272 22894 20324
rect 24026 20272 24032 20324
rect 24084 20312 24090 20324
rect 24765 20315 24823 20321
rect 24765 20312 24777 20315
rect 24084 20284 24777 20312
rect 24084 20272 24090 20284
rect 24765 20281 24777 20284
rect 24811 20281 24823 20315
rect 24765 20275 24823 20281
rect 24857 20315 24915 20321
rect 24857 20281 24869 20315
rect 24903 20281 24915 20315
rect 25056 20312 25084 20343
rect 25314 20340 25320 20392
rect 25372 20380 25378 20392
rect 25593 20383 25651 20389
rect 25593 20380 25605 20383
rect 25372 20352 25605 20380
rect 25372 20340 25378 20352
rect 25593 20349 25605 20352
rect 25639 20349 25651 20383
rect 25774 20380 25780 20392
rect 25735 20352 25780 20380
rect 25593 20343 25651 20349
rect 25774 20340 25780 20352
rect 25832 20340 25838 20392
rect 26418 20380 26424 20392
rect 26379 20352 26424 20380
rect 26418 20340 26424 20352
rect 26476 20340 26482 20392
rect 26602 20340 26608 20392
rect 26660 20340 26666 20392
rect 28442 20380 28448 20392
rect 28403 20352 28448 20380
rect 28442 20340 28448 20352
rect 28500 20340 28506 20392
rect 29549 20383 29607 20389
rect 29549 20349 29561 20383
rect 29595 20349 29607 20383
rect 31312 20380 31340 20547
rect 32030 20544 32036 20596
rect 32088 20584 32094 20596
rect 32125 20587 32183 20593
rect 32125 20584 32137 20587
rect 32088 20556 32137 20584
rect 32088 20544 32094 20556
rect 32125 20553 32137 20556
rect 32171 20553 32183 20587
rect 32125 20547 32183 20553
rect 31757 20383 31815 20389
rect 31757 20380 31769 20383
rect 31312 20352 31769 20380
rect 29549 20343 29607 20349
rect 31757 20349 31769 20352
rect 31803 20349 31815 20383
rect 31757 20343 31815 20349
rect 31941 20383 31999 20389
rect 31941 20349 31953 20383
rect 31987 20380 31999 20383
rect 32214 20380 32220 20392
rect 31987 20352 32220 20380
rect 31987 20349 31999 20352
rect 31941 20343 31999 20349
rect 26620 20312 26648 20340
rect 25056 20284 26648 20312
rect 29564 20312 29592 20343
rect 32214 20340 32220 20352
rect 32272 20340 32278 20392
rect 29822 20312 29828 20324
rect 29564 20284 29828 20312
rect 24857 20275 24915 20281
rect 12986 20244 12992 20256
rect 10336 20216 12992 20244
rect 12986 20204 12992 20216
rect 13044 20204 13050 20256
rect 13449 20247 13507 20253
rect 13449 20213 13461 20247
rect 13495 20244 13507 20247
rect 13906 20244 13912 20256
rect 13495 20216 13912 20244
rect 13495 20213 13507 20216
rect 13449 20207 13507 20213
rect 13906 20204 13912 20216
rect 13964 20204 13970 20256
rect 14090 20244 14096 20256
rect 14051 20216 14096 20244
rect 14090 20204 14096 20216
rect 14148 20204 14154 20256
rect 14826 20204 14832 20256
rect 14884 20244 14890 20256
rect 18414 20244 18420 20256
rect 14884 20216 18420 20244
rect 14884 20204 14890 20216
rect 18414 20204 18420 20216
rect 18472 20204 18478 20256
rect 19058 20204 19064 20256
rect 19116 20244 19122 20256
rect 20162 20244 20168 20256
rect 19116 20216 20168 20244
rect 19116 20204 19122 20216
rect 20162 20204 20168 20216
rect 20220 20204 20226 20256
rect 23566 20204 23572 20256
rect 23624 20244 23630 20256
rect 24489 20247 24547 20253
rect 24489 20244 24501 20247
rect 23624 20216 24501 20244
rect 23624 20204 23630 20216
rect 24489 20213 24501 20216
rect 24535 20213 24547 20247
rect 24872 20244 24900 20275
rect 29822 20272 29828 20284
rect 29880 20272 29886 20324
rect 32582 20312 32588 20324
rect 31050 20284 32588 20312
rect 32582 20272 32588 20284
rect 32640 20272 32646 20324
rect 25590 20244 25596 20256
rect 24872 20216 25596 20244
rect 24489 20207 24547 20213
rect 25590 20204 25596 20216
rect 25648 20204 25654 20256
rect 27614 20204 27620 20256
rect 27672 20244 27678 20256
rect 28537 20247 28595 20253
rect 28537 20244 28549 20247
rect 27672 20216 28549 20244
rect 27672 20204 27678 20216
rect 28537 20213 28549 20216
rect 28583 20213 28595 20247
rect 28537 20207 28595 20213
rect 1104 20154 34316 20176
rect 1104 20102 12052 20154
rect 12104 20102 12116 20154
rect 12168 20102 12180 20154
rect 12232 20102 12244 20154
rect 12296 20102 23123 20154
rect 23175 20102 23187 20154
rect 23239 20102 23251 20154
rect 23303 20102 23315 20154
rect 23367 20102 34316 20154
rect 1104 20080 34316 20102
rect 3050 20040 3056 20052
rect 2963 20012 3056 20040
rect 2976 19981 3004 20012
rect 3050 20000 3056 20012
rect 3108 20040 3114 20052
rect 3326 20040 3332 20052
rect 3108 20012 3332 20040
rect 3108 20000 3114 20012
rect 3326 20000 3332 20012
rect 3384 20000 3390 20052
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 4914 20043 4972 20049
rect 4914 20040 4926 20043
rect 4212 20012 4926 20040
rect 4212 20000 4218 20012
rect 4914 20009 4926 20012
rect 4960 20009 4972 20043
rect 4914 20003 4972 20009
rect 5077 20043 5135 20049
rect 5077 20009 5089 20043
rect 5123 20040 5135 20043
rect 5442 20040 5448 20052
rect 5123 20012 5448 20040
rect 5123 20009 5135 20012
rect 5077 20003 5135 20009
rect 5442 20000 5448 20012
rect 5500 20000 5506 20052
rect 5813 20043 5871 20049
rect 5813 20009 5825 20043
rect 5859 20009 5871 20043
rect 6822 20040 6828 20052
rect 6783 20012 6828 20040
rect 5813 20003 5871 20009
rect 2961 19975 3019 19981
rect 2961 19941 2973 19975
rect 3007 19941 3019 19975
rect 2961 19935 3019 19941
rect 4709 19975 4767 19981
rect 4709 19941 4721 19975
rect 4755 19941 4767 19975
rect 4709 19935 4767 19941
rect 2501 19907 2559 19913
rect 2501 19873 2513 19907
rect 2547 19904 2559 19907
rect 2682 19904 2688 19916
rect 2547 19876 2688 19904
rect 2547 19873 2559 19876
rect 2501 19867 2559 19873
rect 2682 19864 2688 19876
rect 2740 19864 2746 19916
rect 3145 19907 3203 19913
rect 3145 19873 3157 19907
rect 3191 19873 3203 19907
rect 3326 19904 3332 19916
rect 3239 19876 3332 19904
rect 3145 19867 3203 19873
rect 2222 19836 2228 19848
rect 2183 19808 2228 19836
rect 2222 19796 2228 19808
rect 2280 19796 2286 19848
rect 3160 19836 3188 19867
rect 3326 19864 3332 19876
rect 3384 19904 3390 19916
rect 3878 19904 3884 19916
rect 3384 19876 3884 19904
rect 3384 19864 3390 19876
rect 3878 19864 3884 19876
rect 3936 19864 3942 19916
rect 4724 19904 4752 19935
rect 5258 19932 5264 19984
rect 5316 19972 5322 19984
rect 5828 19972 5856 20003
rect 6822 20000 6828 20012
rect 6880 20000 6886 20052
rect 15194 20040 15200 20052
rect 12406 20012 15200 20040
rect 9674 19972 9680 19984
rect 5316 19944 5856 19972
rect 6748 19944 9680 19972
rect 5316 19932 5322 19944
rect 5074 19904 5080 19916
rect 4724 19876 5080 19904
rect 5074 19864 5080 19876
rect 5132 19864 5138 19916
rect 5626 19864 5632 19916
rect 5684 19904 5690 19916
rect 6748 19913 6776 19944
rect 9674 19932 9680 19944
rect 9732 19932 9738 19984
rect 12406 19972 12434 20012
rect 15194 20000 15200 20012
rect 15252 20000 15258 20052
rect 16485 20043 16543 20049
rect 16485 20009 16497 20043
rect 16531 20040 16543 20043
rect 16574 20040 16580 20052
rect 16531 20012 16580 20040
rect 16531 20009 16543 20012
rect 16485 20003 16543 20009
rect 16574 20000 16580 20012
rect 16632 20000 16638 20052
rect 17773 20043 17831 20049
rect 17773 20040 17785 20043
rect 16868 20012 17785 20040
rect 10520 19944 12434 19972
rect 5997 19907 6055 19913
rect 5997 19904 6009 19907
rect 5684 19876 6009 19904
rect 5684 19864 5690 19876
rect 5997 19873 6009 19876
rect 6043 19904 6055 19907
rect 6733 19907 6791 19913
rect 6733 19904 6745 19907
rect 6043 19876 6745 19904
rect 6043 19873 6055 19876
rect 5997 19867 6055 19873
rect 6733 19873 6745 19876
rect 6779 19873 6791 19907
rect 9766 19904 9772 19916
rect 9727 19876 9772 19904
rect 6733 19867 6791 19873
rect 9766 19864 9772 19876
rect 9824 19864 9830 19916
rect 10134 19904 10140 19916
rect 10095 19876 10140 19904
rect 10134 19864 10140 19876
rect 10192 19864 10198 19916
rect 10520 19913 10548 19944
rect 12526 19932 12532 19984
rect 12584 19972 12590 19984
rect 12584 19944 14136 19972
rect 12584 19932 12590 19944
rect 14108 19916 14136 19944
rect 16298 19932 16304 19984
rect 16356 19972 16362 19984
rect 16868 19972 16896 20012
rect 17773 20009 17785 20012
rect 17819 20040 17831 20043
rect 19058 20040 19064 20052
rect 17819 20012 19064 20040
rect 17819 20009 17831 20012
rect 17773 20003 17831 20009
rect 19058 20000 19064 20012
rect 19116 20000 19122 20052
rect 20346 20000 20352 20052
rect 20404 20040 20410 20052
rect 20404 20012 25697 20040
rect 20404 20000 20410 20012
rect 18966 19972 18972 19984
rect 16356 19944 16896 19972
rect 16356 19932 16362 19944
rect 10505 19907 10563 19913
rect 10505 19873 10517 19907
rect 10551 19873 10563 19907
rect 10686 19904 10692 19916
rect 10647 19876 10692 19904
rect 10505 19867 10563 19873
rect 10686 19864 10692 19876
rect 10744 19864 10750 19916
rect 11241 19907 11299 19913
rect 11241 19873 11253 19907
rect 11287 19904 11299 19907
rect 12161 19907 12219 19913
rect 12161 19904 12173 19907
rect 11287 19876 12173 19904
rect 11287 19873 11299 19876
rect 11241 19867 11299 19873
rect 12161 19873 12173 19876
rect 12207 19873 12219 19907
rect 12161 19867 12219 19873
rect 12250 19864 12256 19916
rect 12308 19904 12314 19916
rect 12345 19907 12403 19913
rect 12345 19904 12357 19907
rect 12308 19876 12357 19904
rect 12308 19864 12314 19876
rect 12345 19873 12357 19876
rect 12391 19904 12403 19907
rect 12802 19904 12808 19916
rect 12391 19876 12808 19904
rect 12391 19873 12403 19876
rect 12345 19867 12403 19873
rect 12802 19864 12808 19876
rect 12860 19864 12866 19916
rect 12989 19907 13047 19913
rect 12989 19873 13001 19907
rect 13035 19873 13047 19907
rect 12989 19867 13047 19873
rect 4706 19836 4712 19848
rect 3160 19808 4712 19836
rect 4706 19796 4712 19808
rect 4764 19796 4770 19848
rect 7098 19796 7104 19848
rect 7156 19836 7162 19848
rect 10229 19839 10287 19845
rect 10229 19836 10241 19839
rect 7156 19808 10241 19836
rect 7156 19796 7162 19808
rect 10229 19805 10241 19808
rect 10275 19805 10287 19839
rect 10229 19799 10287 19805
rect 11790 19796 11796 19848
rect 11848 19836 11854 19848
rect 13004 19836 13032 19867
rect 14090 19864 14096 19916
rect 14148 19904 14154 19916
rect 14737 19907 14795 19913
rect 14737 19904 14749 19907
rect 14148 19876 14749 19904
rect 14148 19864 14154 19876
rect 14737 19873 14749 19876
rect 14783 19873 14795 19907
rect 14737 19867 14795 19873
rect 14921 19907 14979 19913
rect 14921 19873 14933 19907
rect 14967 19873 14979 19907
rect 14921 19867 14979 19873
rect 11848 19808 13032 19836
rect 11848 19796 11854 19808
rect 1946 19728 1952 19780
rect 2004 19768 2010 19780
rect 2004 19740 12434 19768
rect 2004 19728 2010 19740
rect 1670 19660 1676 19712
rect 1728 19700 1734 19712
rect 2317 19703 2375 19709
rect 2317 19700 2329 19703
rect 1728 19672 2329 19700
rect 1728 19660 1734 19672
rect 2317 19669 2329 19672
rect 2363 19669 2375 19703
rect 2317 19663 2375 19669
rect 2409 19703 2467 19709
rect 2409 19669 2421 19703
rect 2455 19700 2467 19703
rect 3142 19700 3148 19712
rect 2455 19672 3148 19700
rect 2455 19669 2467 19672
rect 2409 19663 2467 19669
rect 3142 19660 3148 19672
rect 3200 19660 3206 19712
rect 4062 19660 4068 19712
rect 4120 19700 4126 19712
rect 4893 19703 4951 19709
rect 4893 19700 4905 19703
rect 4120 19672 4905 19700
rect 4120 19660 4126 19672
rect 4893 19669 4905 19672
rect 4939 19669 4951 19703
rect 12406 19700 12434 19740
rect 12894 19728 12900 19780
rect 12952 19768 12958 19780
rect 13173 19771 13231 19777
rect 13173 19768 13185 19771
rect 12952 19740 13185 19768
rect 12952 19728 12958 19740
rect 13173 19737 13185 19740
rect 13219 19768 13231 19771
rect 14936 19768 14964 19867
rect 15010 19864 15016 19916
rect 15068 19904 15074 19916
rect 15151 19907 15209 19913
rect 15068 19876 15113 19904
rect 15068 19864 15074 19876
rect 15151 19873 15163 19907
rect 15197 19904 15209 19907
rect 16025 19907 16083 19913
rect 15197 19876 15332 19904
rect 15197 19873 15209 19876
rect 15151 19867 15209 19873
rect 15304 19836 15332 19876
rect 16025 19873 16037 19907
rect 16071 19904 16083 19907
rect 16758 19904 16764 19916
rect 16071 19876 16764 19904
rect 16071 19873 16083 19876
rect 16025 19867 16083 19873
rect 16758 19864 16764 19876
rect 16816 19864 16822 19916
rect 16868 19913 16896 19944
rect 17144 19944 18972 19972
rect 17144 19913 17172 19944
rect 18966 19932 18972 19944
rect 19024 19932 19030 19984
rect 21358 19932 21364 19984
rect 21416 19932 21422 19984
rect 24213 19975 24271 19981
rect 24213 19941 24225 19975
rect 24259 19972 24271 19975
rect 25314 19972 25320 19984
rect 24259 19944 25320 19972
rect 24259 19941 24271 19944
rect 24213 19935 24271 19941
rect 25314 19932 25320 19944
rect 25372 19972 25378 19984
rect 25669 19972 25697 20012
rect 26510 20000 26516 20052
rect 26568 20040 26574 20052
rect 26568 20012 26613 20040
rect 26568 20000 26574 20012
rect 27065 19975 27123 19981
rect 25372 19932 25381 19972
rect 25669 19944 25912 19972
rect 16853 19907 16911 19913
rect 16853 19873 16865 19907
rect 16899 19873 16911 19907
rect 16853 19867 16911 19873
rect 16945 19907 17003 19913
rect 16945 19873 16957 19907
rect 16991 19873 17003 19907
rect 16945 19867 17003 19873
rect 17129 19907 17187 19913
rect 17129 19873 17141 19907
rect 17175 19873 17187 19907
rect 17129 19867 17187 19873
rect 13219 19740 14964 19768
rect 15028 19808 15332 19836
rect 13219 19737 13231 19740
rect 13173 19731 13231 19737
rect 14826 19700 14832 19712
rect 12406 19672 14832 19700
rect 4893 19663 4951 19669
rect 14826 19660 14832 19672
rect 14884 19660 14890 19712
rect 14918 19660 14924 19712
rect 14976 19700 14982 19712
rect 15028 19700 15056 19808
rect 16114 19728 16120 19780
rect 16172 19768 16178 19780
rect 16960 19768 16988 19867
rect 17310 19864 17316 19916
rect 17368 19904 17374 19916
rect 17589 19907 17647 19913
rect 17589 19904 17601 19907
rect 17368 19876 17601 19904
rect 17368 19864 17374 19876
rect 17589 19873 17601 19876
rect 17635 19873 17647 19907
rect 17589 19867 17647 19873
rect 17862 19864 17868 19916
rect 17920 19904 17926 19916
rect 22741 19907 22799 19913
rect 17920 19876 17965 19904
rect 17920 19864 17926 19876
rect 22741 19873 22753 19907
rect 22787 19873 22799 19907
rect 22741 19867 22799 19873
rect 22925 19907 22983 19913
rect 22925 19873 22937 19907
rect 22971 19904 22983 19907
rect 23014 19904 23020 19916
rect 22971 19876 23020 19904
rect 22971 19873 22983 19876
rect 22925 19867 22983 19873
rect 20254 19796 20260 19848
rect 20312 19836 20318 19848
rect 20349 19839 20407 19845
rect 20349 19836 20361 19839
rect 20312 19808 20361 19836
rect 20312 19796 20318 19808
rect 20349 19805 20361 19808
rect 20395 19805 20407 19839
rect 20349 19799 20407 19805
rect 20625 19839 20683 19845
rect 20625 19805 20637 19839
rect 20671 19836 20683 19839
rect 20714 19836 20720 19848
rect 20671 19808 20720 19836
rect 20671 19805 20683 19808
rect 20625 19799 20683 19805
rect 20714 19796 20720 19808
rect 20772 19796 20778 19848
rect 22756 19836 22784 19867
rect 23014 19864 23020 19876
rect 23072 19864 23078 19916
rect 24302 19904 24308 19916
rect 24263 19876 24308 19904
rect 24302 19864 24308 19876
rect 24360 19864 24366 19916
rect 24762 19864 24768 19916
rect 24820 19904 24826 19916
rect 25353 19913 25381 19932
rect 25225 19907 25283 19913
rect 25225 19904 25237 19907
rect 24820 19876 25237 19904
rect 24820 19864 24826 19876
rect 25225 19873 25237 19876
rect 25271 19873 25283 19907
rect 25353 19907 25421 19913
rect 25353 19876 25375 19907
rect 25225 19867 25283 19873
rect 25363 19873 25375 19876
rect 25409 19873 25421 19907
rect 25363 19867 25421 19873
rect 25593 19907 25651 19913
rect 25593 19873 25605 19907
rect 25639 19904 25651 19907
rect 25774 19904 25780 19916
rect 25639 19876 25780 19904
rect 25639 19873 25651 19876
rect 25593 19867 25651 19873
rect 25774 19864 25780 19876
rect 25832 19864 25838 19916
rect 25884 19904 25912 19944
rect 27065 19941 27077 19975
rect 27111 19972 27123 19975
rect 27614 19972 27620 19984
rect 27111 19944 27620 19972
rect 27111 19941 27123 19944
rect 27065 19935 27123 19941
rect 27614 19932 27620 19944
rect 27672 19932 27678 19984
rect 32582 19932 32588 19984
rect 32640 19932 32646 19984
rect 26418 19904 26424 19916
rect 25884 19876 26424 19904
rect 26418 19864 26424 19876
rect 26476 19864 26482 19916
rect 27246 19904 27252 19916
rect 27207 19876 27252 19904
rect 27246 19864 27252 19876
rect 27304 19864 27310 19916
rect 27338 19864 27344 19916
rect 27396 19904 27402 19916
rect 27433 19907 27491 19913
rect 27433 19904 27445 19907
rect 27396 19876 27445 19904
rect 27396 19864 27402 19876
rect 27433 19873 27445 19876
rect 27479 19904 27491 19907
rect 28537 19907 28595 19913
rect 28537 19904 28549 19907
rect 27479 19876 28549 19904
rect 27479 19873 27491 19876
rect 27433 19867 27491 19873
rect 28537 19873 28549 19876
rect 28583 19873 28595 19907
rect 28537 19867 28595 19873
rect 25682 19836 25688 19848
rect 22756 19808 25688 19836
rect 18690 19768 18696 19780
rect 16172 19740 18696 19768
rect 16172 19728 16178 19740
rect 18690 19728 18696 19740
rect 18748 19728 18754 19780
rect 21634 19728 21640 19780
rect 21692 19768 21698 19780
rect 22756 19768 22784 19808
rect 25682 19796 25688 19808
rect 25740 19796 25746 19848
rect 26436 19836 26464 19864
rect 28258 19836 28264 19848
rect 26436 19808 28264 19836
rect 28258 19796 28264 19808
rect 28316 19796 28322 19848
rect 28442 19836 28448 19848
rect 28403 19808 28448 19836
rect 28442 19796 28448 19808
rect 28500 19796 28506 19848
rect 31754 19796 31760 19848
rect 31812 19836 31818 19848
rect 31849 19839 31907 19845
rect 31849 19836 31861 19839
rect 31812 19808 31861 19836
rect 31812 19796 31818 19808
rect 31849 19805 31861 19808
rect 31895 19805 31907 19839
rect 32122 19836 32128 19848
rect 32083 19808 32128 19836
rect 31849 19799 31907 19805
rect 32122 19796 32128 19808
rect 32180 19796 32186 19848
rect 21692 19740 22784 19768
rect 21692 19728 21698 19740
rect 14976 19672 15056 19700
rect 15381 19703 15439 19709
rect 14976 19660 14982 19672
rect 15381 19669 15393 19703
rect 15427 19700 15439 19703
rect 15746 19700 15752 19712
rect 15427 19672 15752 19700
rect 15427 19669 15439 19672
rect 15381 19663 15439 19669
rect 15746 19660 15752 19672
rect 15804 19660 15810 19712
rect 15933 19703 15991 19709
rect 15933 19669 15945 19703
rect 15979 19700 15991 19703
rect 16022 19700 16028 19712
rect 15979 19672 16028 19700
rect 15979 19669 15991 19672
rect 15933 19663 15991 19669
rect 16022 19660 16028 19672
rect 16080 19660 16086 19712
rect 16574 19660 16580 19712
rect 16632 19700 16638 19712
rect 17589 19703 17647 19709
rect 17589 19700 17601 19703
rect 16632 19672 17601 19700
rect 16632 19660 16638 19672
rect 17589 19669 17601 19672
rect 17635 19669 17647 19703
rect 17589 19663 17647 19669
rect 22094 19660 22100 19712
rect 22152 19700 22158 19712
rect 22152 19672 22197 19700
rect 22152 19660 22158 19672
rect 22646 19660 22652 19712
rect 22704 19700 22710 19712
rect 22741 19703 22799 19709
rect 22741 19700 22753 19703
rect 22704 19672 22753 19700
rect 22704 19660 22710 19672
rect 22741 19669 22753 19672
rect 22787 19669 22799 19703
rect 22741 19663 22799 19669
rect 28905 19703 28963 19709
rect 28905 19669 28917 19703
rect 28951 19700 28963 19703
rect 29546 19700 29552 19712
rect 28951 19672 29552 19700
rect 28951 19669 28963 19672
rect 28905 19663 28963 19669
rect 29546 19660 29552 19672
rect 29604 19660 29610 19712
rect 33594 19700 33600 19712
rect 33555 19672 33600 19700
rect 33594 19660 33600 19672
rect 33652 19660 33658 19712
rect 1104 19610 34316 19632
rect 1104 19558 6517 19610
rect 6569 19558 6581 19610
rect 6633 19558 6645 19610
rect 6697 19558 6709 19610
rect 6761 19558 17588 19610
rect 17640 19558 17652 19610
rect 17704 19558 17716 19610
rect 17768 19558 17780 19610
rect 17832 19558 28658 19610
rect 28710 19558 28722 19610
rect 28774 19558 28786 19610
rect 28838 19558 28850 19610
rect 28902 19558 34316 19610
rect 1104 19536 34316 19558
rect 3145 19499 3203 19505
rect 3145 19465 3157 19499
rect 3191 19496 3203 19499
rect 3326 19496 3332 19508
rect 3191 19468 3332 19496
rect 3191 19465 3203 19468
rect 3145 19459 3203 19465
rect 3326 19456 3332 19468
rect 3384 19456 3390 19508
rect 3970 19496 3976 19508
rect 3931 19468 3976 19496
rect 3970 19456 3976 19468
rect 4028 19456 4034 19508
rect 4430 19456 4436 19508
rect 4488 19496 4494 19508
rect 4525 19499 4583 19505
rect 4525 19496 4537 19499
rect 4488 19468 4537 19496
rect 4488 19456 4494 19468
rect 4525 19465 4537 19468
rect 4571 19465 4583 19499
rect 4525 19459 4583 19465
rect 10502 19456 10508 19508
rect 10560 19496 10566 19508
rect 12250 19496 12256 19508
rect 10560 19468 10824 19496
rect 12211 19468 12256 19496
rect 10560 19456 10566 19468
rect 9953 19431 10011 19437
rect 9953 19397 9965 19431
rect 9999 19428 10011 19431
rect 10686 19428 10692 19440
rect 9999 19400 10692 19428
rect 9999 19397 10011 19400
rect 9953 19391 10011 19397
rect 10686 19388 10692 19400
rect 10744 19388 10750 19440
rect 10796 19428 10824 19468
rect 12250 19456 12256 19468
rect 12308 19456 12314 19508
rect 13170 19496 13176 19508
rect 13131 19468 13176 19496
rect 13170 19456 13176 19468
rect 13228 19456 13234 19508
rect 13538 19496 13544 19508
rect 13499 19468 13544 19496
rect 13538 19456 13544 19468
rect 13596 19456 13602 19508
rect 14826 19456 14832 19508
rect 14884 19496 14890 19508
rect 15838 19496 15844 19508
rect 14884 19468 15844 19496
rect 14884 19456 14890 19468
rect 15838 19456 15844 19468
rect 15896 19496 15902 19508
rect 17773 19499 17831 19505
rect 17773 19496 17785 19499
rect 15896 19468 17785 19496
rect 15896 19456 15902 19468
rect 17773 19465 17785 19468
rect 17819 19496 17831 19499
rect 21634 19496 21640 19508
rect 17819 19468 21640 19496
rect 17819 19465 17831 19468
rect 17773 19459 17831 19465
rect 21634 19456 21640 19468
rect 21692 19456 21698 19508
rect 24302 19456 24308 19508
rect 24360 19496 24366 19508
rect 25041 19499 25099 19505
rect 25041 19496 25053 19499
rect 24360 19468 25053 19496
rect 24360 19456 24366 19468
rect 25041 19465 25053 19468
rect 25087 19496 25099 19499
rect 27246 19496 27252 19508
rect 25087 19468 27252 19496
rect 25087 19465 25099 19468
rect 25041 19459 25099 19465
rect 27246 19456 27252 19468
rect 27304 19456 27310 19508
rect 13814 19428 13820 19440
rect 10796 19400 13820 19428
rect 13814 19388 13820 19400
rect 13872 19388 13878 19440
rect 14642 19388 14648 19440
rect 14700 19428 14706 19440
rect 14921 19431 14979 19437
rect 14921 19428 14933 19431
rect 14700 19400 14933 19428
rect 14700 19388 14706 19400
rect 14921 19397 14933 19400
rect 14967 19397 14979 19431
rect 14921 19391 14979 19397
rect 15059 19431 15117 19437
rect 15059 19397 15071 19431
rect 15105 19428 15117 19431
rect 16022 19428 16028 19440
rect 15105 19400 16028 19428
rect 15105 19397 15117 19400
rect 15059 19391 15117 19397
rect 16022 19388 16028 19400
rect 16080 19388 16086 19440
rect 32214 19388 32220 19440
rect 32272 19428 32278 19440
rect 33137 19431 33195 19437
rect 33137 19428 33149 19431
rect 32272 19400 33149 19428
rect 32272 19388 32278 19400
rect 33137 19397 33149 19400
rect 33183 19397 33195 19431
rect 33137 19391 33195 19397
rect 1670 19360 1676 19372
rect 1631 19332 1676 19360
rect 1670 19320 1676 19332
rect 1728 19320 1734 19372
rect 5626 19360 5632 19372
rect 5587 19332 5632 19360
rect 5626 19320 5632 19332
rect 5684 19320 5690 19372
rect 7098 19360 7104 19372
rect 7059 19332 7104 19360
rect 7098 19320 7104 19332
rect 7156 19320 7162 19372
rect 12894 19360 12900 19372
rect 9692 19332 10640 19360
rect 1394 19292 1400 19304
rect 1307 19264 1400 19292
rect 1394 19252 1400 19264
rect 1452 19252 1458 19304
rect 4522 19292 4528 19304
rect 3620 19264 3832 19292
rect 4483 19264 4528 19292
rect 1412 19224 1440 19252
rect 1412 19196 1532 19224
rect 1504 19156 1532 19196
rect 2406 19184 2412 19236
rect 2464 19184 2470 19236
rect 3620 19156 3648 19264
rect 3697 19227 3755 19233
rect 3697 19193 3709 19227
rect 3743 19193 3755 19227
rect 3804 19224 3832 19264
rect 4522 19252 4528 19264
rect 4580 19252 4586 19304
rect 4706 19292 4712 19304
rect 4667 19264 4712 19292
rect 4706 19252 4712 19264
rect 4764 19252 4770 19304
rect 4801 19295 4859 19301
rect 4801 19261 4813 19295
rect 4847 19261 4859 19295
rect 4801 19255 4859 19261
rect 4816 19224 4844 19255
rect 5074 19252 5080 19304
rect 5132 19292 5138 19304
rect 5261 19295 5319 19301
rect 5261 19292 5273 19295
rect 5132 19264 5273 19292
rect 5132 19252 5138 19264
rect 5261 19261 5273 19264
rect 5307 19261 5319 19295
rect 5534 19292 5540 19304
rect 5495 19264 5540 19292
rect 5261 19255 5319 19261
rect 5534 19252 5540 19264
rect 5592 19252 5598 19304
rect 6825 19295 6883 19301
rect 6825 19261 6837 19295
rect 6871 19261 6883 19295
rect 6825 19255 6883 19261
rect 5552 19224 5580 19252
rect 3804 19196 4752 19224
rect 4816 19196 5580 19224
rect 3697 19187 3755 19193
rect 1504 19128 3648 19156
rect 3712 19156 3740 19187
rect 4154 19156 4160 19168
rect 3712 19128 4160 19156
rect 4154 19116 4160 19128
rect 4212 19116 4218 19168
rect 4724 19156 4752 19196
rect 6840 19156 6868 19255
rect 8938 19252 8944 19304
rect 8996 19292 9002 19304
rect 9033 19295 9091 19301
rect 9033 19292 9045 19295
rect 8996 19264 9045 19292
rect 8996 19252 9002 19264
rect 9033 19261 9045 19264
rect 9079 19261 9091 19295
rect 9033 19255 9091 19261
rect 9217 19295 9275 19301
rect 9217 19261 9229 19295
rect 9263 19292 9275 19295
rect 9306 19292 9312 19304
rect 9263 19264 9312 19292
rect 9263 19261 9275 19264
rect 9217 19255 9275 19261
rect 9306 19252 9312 19264
rect 9364 19252 9370 19304
rect 9582 19292 9588 19304
rect 9543 19264 9588 19292
rect 9582 19252 9588 19264
rect 9640 19292 9646 19304
rect 9692 19292 9720 19332
rect 9640 19264 9720 19292
rect 9769 19295 9827 19301
rect 9640 19252 9646 19264
rect 9769 19261 9781 19295
rect 9815 19261 9827 19295
rect 10042 19292 10048 19304
rect 10003 19264 10048 19292
rect 9769 19255 9827 19261
rect 7006 19184 7012 19236
rect 7064 19224 7070 19236
rect 7064 19210 7590 19224
rect 7064 19196 7604 19210
rect 7064 19184 7070 19196
rect 4724 19128 6868 19156
rect 7576 19156 7604 19196
rect 8386 19156 8392 19168
rect 7576 19128 8392 19156
rect 8386 19116 8392 19128
rect 8444 19116 8450 19168
rect 8478 19116 8484 19168
rect 8536 19156 8542 19168
rect 8573 19159 8631 19165
rect 8573 19156 8585 19159
rect 8536 19128 8585 19156
rect 8536 19116 8542 19128
rect 8573 19125 8585 19128
rect 8619 19156 8631 19159
rect 9784 19156 9812 19255
rect 10042 19252 10048 19264
rect 10100 19252 10106 19304
rect 10612 19301 10640 19332
rect 12360 19332 12900 19360
rect 10505 19295 10563 19301
rect 10505 19261 10517 19295
rect 10551 19261 10563 19295
rect 10505 19255 10563 19261
rect 10597 19295 10655 19301
rect 10597 19261 10609 19295
rect 10643 19261 10655 19295
rect 10597 19255 10655 19261
rect 9858 19184 9864 19236
rect 9916 19224 9922 19236
rect 10520 19224 10548 19255
rect 11790 19252 11796 19304
rect 11848 19292 11854 19304
rect 12161 19295 12219 19301
rect 12161 19292 12173 19295
rect 11848 19264 12173 19292
rect 11848 19252 11854 19264
rect 12161 19261 12173 19264
rect 12207 19261 12219 19295
rect 12161 19255 12219 19261
rect 9916 19196 10548 19224
rect 9916 19184 9922 19196
rect 11514 19184 11520 19236
rect 11572 19224 11578 19236
rect 12360 19224 12388 19332
rect 12894 19320 12900 19332
rect 12952 19320 12958 19372
rect 13630 19320 13636 19372
rect 13688 19360 13694 19372
rect 14829 19363 14887 19369
rect 14829 19360 14841 19363
rect 13688 19332 14841 19360
rect 13688 19320 13694 19332
rect 14829 19329 14841 19332
rect 14875 19329 14887 19363
rect 15381 19363 15439 19369
rect 15381 19360 15393 19363
rect 14829 19323 14887 19329
rect 15304 19332 15393 19360
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19261 12495 19295
rect 13354 19292 13360 19304
rect 13315 19264 13360 19292
rect 12437 19255 12495 19261
rect 11572 19196 12388 19224
rect 11572 19184 11578 19196
rect 8619 19128 9812 19156
rect 8619 19125 8631 19128
rect 8573 19119 8631 19125
rect 10686 19116 10692 19168
rect 10744 19156 10750 19168
rect 12452 19156 12480 19255
rect 13354 19252 13360 19264
rect 13412 19252 13418 19304
rect 13446 19252 13452 19304
rect 13504 19292 13510 19304
rect 13541 19295 13599 19301
rect 13541 19292 13553 19295
rect 13504 19264 13553 19292
rect 13504 19252 13510 19264
rect 13541 19261 13553 19264
rect 13587 19261 13599 19295
rect 13541 19255 13599 19261
rect 13906 19252 13912 19304
rect 13964 19292 13970 19304
rect 15304 19292 15332 19332
rect 15381 19329 15393 19332
rect 15427 19329 15439 19363
rect 15381 19323 15439 19329
rect 15746 19320 15752 19372
rect 15804 19360 15810 19372
rect 16393 19363 16451 19369
rect 16393 19360 16405 19363
rect 15804 19332 16405 19360
rect 15804 19320 15810 19332
rect 16393 19329 16405 19332
rect 16439 19329 16451 19363
rect 16393 19323 16451 19329
rect 20622 19320 20628 19372
rect 20680 19360 20686 19372
rect 20717 19363 20775 19369
rect 20717 19360 20729 19363
rect 20680 19332 20729 19360
rect 20680 19320 20686 19332
rect 20717 19329 20729 19332
rect 20763 19329 20775 19363
rect 20717 19323 20775 19329
rect 15470 19292 15476 19304
rect 13964 19264 15332 19292
rect 15431 19264 15476 19292
rect 13964 19252 13970 19264
rect 15470 19252 15476 19264
rect 15528 19252 15534 19304
rect 15838 19292 15844 19304
rect 15799 19264 15844 19292
rect 15838 19252 15844 19264
rect 15896 19252 15902 19304
rect 16114 19292 16120 19304
rect 16075 19264 16120 19292
rect 16114 19252 16120 19264
rect 16172 19252 16178 19304
rect 16301 19295 16359 19301
rect 16301 19261 16313 19295
rect 16347 19261 16359 19295
rect 19886 19292 19892 19304
rect 19847 19264 19892 19292
rect 16301 19255 16359 19261
rect 13998 19184 14004 19236
rect 14056 19224 14062 19236
rect 14461 19227 14519 19233
rect 14461 19224 14473 19227
rect 14056 19196 14473 19224
rect 14056 19184 14062 19196
rect 14461 19193 14473 19196
rect 14507 19193 14519 19227
rect 14461 19187 14519 19193
rect 15010 19184 15016 19236
rect 15068 19224 15074 19236
rect 15197 19227 15255 19233
rect 15197 19224 15209 19227
rect 15068 19196 15209 19224
rect 15068 19184 15074 19196
rect 15197 19193 15209 19196
rect 15243 19193 15255 19227
rect 15197 19187 15255 19193
rect 15286 19184 15292 19236
rect 15344 19224 15350 19236
rect 15565 19227 15623 19233
rect 15344 19196 15389 19224
rect 15344 19184 15350 19196
rect 15565 19193 15577 19227
rect 15611 19193 15623 19227
rect 15565 19187 15623 19193
rect 15657 19227 15715 19233
rect 15657 19193 15669 19227
rect 15703 19224 15715 19227
rect 15746 19224 15752 19236
rect 15703 19196 15752 19224
rect 15703 19193 15715 19196
rect 15657 19187 15715 19193
rect 14826 19156 14832 19168
rect 10744 19128 14832 19156
rect 10744 19116 10750 19128
rect 14826 19116 14832 19128
rect 14884 19116 14890 19168
rect 15102 19116 15108 19168
rect 15160 19156 15166 19168
rect 15580 19156 15608 19187
rect 15746 19184 15752 19196
rect 15804 19184 15810 19236
rect 16316 19224 16344 19255
rect 19886 19252 19892 19264
rect 19944 19252 19950 19304
rect 20165 19295 20223 19301
rect 20165 19261 20177 19295
rect 20211 19292 20223 19295
rect 20346 19292 20352 19304
rect 20211 19264 20352 19292
rect 20211 19261 20223 19264
rect 20165 19255 20223 19261
rect 20346 19252 20352 19264
rect 20404 19252 20410 19304
rect 20806 19294 20812 19346
rect 20864 19294 20870 19346
rect 20898 19320 20904 19372
rect 20956 19360 20962 19372
rect 20956 19332 21001 19360
rect 20956 19320 20962 19332
rect 22462 19320 22468 19372
rect 22520 19360 22526 19372
rect 22833 19363 22891 19369
rect 22833 19360 22845 19363
rect 22520 19332 22845 19360
rect 22520 19320 22526 19332
rect 22833 19329 22845 19332
rect 22879 19329 22891 19363
rect 23566 19360 23572 19372
rect 23527 19332 23572 19360
rect 22833 19323 22891 19329
rect 23566 19320 23572 19332
rect 23624 19320 23630 19372
rect 30834 19320 30840 19372
rect 30892 19360 30898 19372
rect 31021 19363 31079 19369
rect 31021 19360 31033 19363
rect 30892 19332 31033 19360
rect 30892 19320 30898 19332
rect 31021 19329 31033 19332
rect 31067 19329 31079 19363
rect 31202 19360 31208 19372
rect 31163 19332 31208 19360
rect 31021 19323 31079 19329
rect 31202 19320 31208 19332
rect 31260 19320 31266 19372
rect 33505 19363 33563 19369
rect 33505 19329 33517 19363
rect 33551 19360 33563 19363
rect 33594 19360 33600 19372
rect 33551 19332 33600 19360
rect 33551 19329 33563 19332
rect 33505 19323 33563 19329
rect 33594 19320 33600 19332
rect 33652 19320 33658 19372
rect 16574 19224 16580 19236
rect 16316 19196 16580 19224
rect 16574 19184 16580 19196
rect 16632 19184 16638 19236
rect 17770 19184 17776 19236
rect 17828 19224 17834 19236
rect 18049 19227 18107 19233
rect 18049 19224 18061 19227
rect 17828 19196 18061 19224
rect 17828 19184 17834 19196
rect 18049 19193 18061 19196
rect 18095 19193 18107 19227
rect 20714 19224 20720 19236
rect 20675 19196 20720 19224
rect 18049 19187 18107 19193
rect 20714 19184 20720 19196
rect 20772 19184 20778 19236
rect 20824 19224 20852 19294
rect 20990 19292 20996 19304
rect 20951 19264 20996 19292
rect 20990 19252 20996 19264
rect 21048 19292 21054 19304
rect 21545 19295 21603 19301
rect 21545 19292 21557 19295
rect 21048 19264 21557 19292
rect 21048 19252 21054 19264
rect 21545 19261 21557 19264
rect 21591 19261 21603 19295
rect 21545 19255 21603 19261
rect 21637 19295 21695 19301
rect 21637 19261 21649 19295
rect 21683 19292 21695 19295
rect 22094 19292 22100 19304
rect 21683 19264 22100 19292
rect 21683 19261 21695 19264
rect 21637 19255 21695 19261
rect 22094 19252 22100 19264
rect 22152 19252 22158 19304
rect 22646 19292 22652 19304
rect 22607 19264 22652 19292
rect 22646 19252 22652 19264
rect 22704 19252 22710 19304
rect 22738 19252 22744 19304
rect 22796 19292 22802 19304
rect 23293 19295 23351 19301
rect 23293 19292 23305 19295
rect 22796 19264 23305 19292
rect 22796 19252 22802 19264
rect 23293 19261 23305 19264
rect 23339 19261 23351 19295
rect 23293 19255 23351 19261
rect 25314 19252 25320 19304
rect 25372 19292 25378 19304
rect 25593 19295 25651 19301
rect 25593 19292 25605 19295
rect 25372 19264 25605 19292
rect 25372 19252 25378 19264
rect 25593 19261 25605 19264
rect 25639 19261 25651 19295
rect 25593 19255 25651 19261
rect 26513 19295 26571 19301
rect 26513 19261 26525 19295
rect 26559 19261 26571 19295
rect 26513 19255 26571 19261
rect 22554 19224 22560 19236
rect 20824 19196 22560 19224
rect 22554 19184 22560 19196
rect 22612 19184 22618 19236
rect 22664 19224 22692 19252
rect 23014 19224 23020 19236
rect 22664 19196 23020 19224
rect 23014 19184 23020 19196
rect 23072 19184 23078 19236
rect 23658 19184 23664 19236
rect 23716 19224 23722 19236
rect 23716 19196 24058 19224
rect 23716 19184 23722 19196
rect 25130 19184 25136 19236
rect 25188 19224 25194 19236
rect 26528 19224 26556 19255
rect 26602 19252 26608 19304
rect 26660 19292 26666 19304
rect 26789 19295 26847 19301
rect 26660 19264 26705 19292
rect 26660 19252 26666 19264
rect 26789 19261 26801 19295
rect 26835 19292 26847 19295
rect 27338 19292 27344 19304
rect 26835 19264 27344 19292
rect 26835 19261 26847 19264
rect 26789 19255 26847 19261
rect 27338 19252 27344 19264
rect 27396 19252 27402 19304
rect 29546 19252 29552 19304
rect 29604 19301 29610 19304
rect 29604 19292 29616 19301
rect 29822 19292 29828 19304
rect 29604 19264 29649 19292
rect 29783 19264 29828 19292
rect 29604 19255 29616 19264
rect 29604 19252 29610 19255
rect 29822 19252 29828 19264
rect 29880 19292 29886 19304
rect 31754 19292 31760 19304
rect 29880 19264 31760 19292
rect 29880 19252 29886 19264
rect 31754 19252 31760 19264
rect 31812 19252 31818 19304
rect 26970 19224 26976 19236
rect 25188 19196 26976 19224
rect 25188 19184 25194 19196
rect 26970 19184 26976 19196
rect 27028 19184 27034 19236
rect 30929 19227 30987 19233
rect 30929 19193 30941 19227
rect 30975 19224 30987 19227
rect 30975 19196 31754 19224
rect 30975 19193 30987 19196
rect 30929 19187 30987 19193
rect 15160 19128 15608 19156
rect 15160 19116 15166 19128
rect 15930 19116 15936 19168
rect 15988 19156 15994 19168
rect 15988 19128 16033 19156
rect 15988 19116 15994 19128
rect 19794 19116 19800 19168
rect 19852 19156 19858 19168
rect 20073 19159 20131 19165
rect 20073 19156 20085 19159
rect 19852 19128 20085 19156
rect 19852 19116 19858 19128
rect 20073 19125 20085 19128
rect 20119 19156 20131 19159
rect 20438 19156 20444 19168
rect 20119 19128 20444 19156
rect 20119 19125 20131 19128
rect 20073 19119 20131 19125
rect 20438 19116 20444 19128
rect 20496 19116 20502 19168
rect 25222 19116 25228 19168
rect 25280 19156 25286 19168
rect 25682 19156 25688 19168
rect 25280 19128 25688 19156
rect 25280 19116 25286 19128
rect 25682 19116 25688 19128
rect 25740 19116 25746 19168
rect 26234 19116 26240 19168
rect 26292 19156 26298 19168
rect 26513 19159 26571 19165
rect 26513 19156 26525 19159
rect 26292 19128 26525 19156
rect 26292 19116 26298 19128
rect 26513 19125 26525 19128
rect 26559 19125 26571 19159
rect 28442 19156 28448 19168
rect 28403 19128 28448 19156
rect 26513 19119 26571 19125
rect 28442 19116 28448 19128
rect 28500 19116 28506 19168
rect 30561 19159 30619 19165
rect 30561 19125 30573 19159
rect 30607 19156 30619 19159
rect 30742 19156 30748 19168
rect 30607 19128 30748 19156
rect 30607 19125 30619 19128
rect 30561 19119 30619 19125
rect 30742 19116 30748 19128
rect 30800 19116 30806 19168
rect 31726 19156 31754 19196
rect 32214 19156 32220 19168
rect 31726 19128 32220 19156
rect 32214 19116 32220 19128
rect 32272 19116 32278 19168
rect 33042 19156 33048 19168
rect 33003 19128 33048 19156
rect 33042 19116 33048 19128
rect 33100 19116 33106 19168
rect 1104 19066 34316 19088
rect 1104 19014 12052 19066
rect 12104 19014 12116 19066
rect 12168 19014 12180 19066
rect 12232 19014 12244 19066
rect 12296 19014 23123 19066
rect 23175 19014 23187 19066
rect 23239 19014 23251 19066
rect 23303 19014 23315 19066
rect 23367 19014 34316 19066
rect 1104 18992 34316 19014
rect 2222 18912 2228 18964
rect 2280 18952 2286 18964
rect 2409 18955 2467 18961
rect 2409 18952 2421 18955
rect 2280 18924 2421 18952
rect 2280 18912 2286 18924
rect 2409 18921 2421 18924
rect 2455 18921 2467 18955
rect 2409 18915 2467 18921
rect 4522 18912 4528 18964
rect 4580 18952 4586 18964
rect 4709 18955 4767 18961
rect 4709 18952 4721 18955
rect 4580 18924 4721 18952
rect 4580 18912 4586 18924
rect 4709 18921 4721 18924
rect 4755 18921 4767 18955
rect 4709 18915 4767 18921
rect 5534 18912 5540 18964
rect 5592 18952 5598 18964
rect 5629 18955 5687 18961
rect 5629 18952 5641 18955
rect 5592 18924 5641 18952
rect 5592 18912 5598 18924
rect 5629 18921 5641 18924
rect 5675 18921 5687 18955
rect 5629 18915 5687 18921
rect 9769 18955 9827 18961
rect 9769 18921 9781 18955
rect 9815 18952 9827 18955
rect 9858 18952 9864 18964
rect 9815 18924 9864 18952
rect 9815 18921 9827 18924
rect 9769 18915 9827 18921
rect 9858 18912 9864 18924
rect 9916 18912 9922 18964
rect 10042 18912 10048 18964
rect 10100 18952 10106 18964
rect 11425 18955 11483 18961
rect 10100 18924 11284 18952
rect 10100 18912 10106 18924
rect 2682 18884 2688 18896
rect 2424 18856 2688 18884
rect 2424 18825 2452 18856
rect 2682 18844 2688 18856
rect 2740 18844 2746 18896
rect 4154 18844 4160 18896
rect 4212 18884 4218 18896
rect 4861 18887 4919 18893
rect 4861 18884 4873 18887
rect 4212 18856 4873 18884
rect 4212 18844 4218 18856
rect 4861 18853 4873 18856
rect 4907 18884 4919 18887
rect 5074 18884 5080 18896
rect 4907 18853 4936 18884
rect 5035 18856 5080 18884
rect 4861 18847 4936 18853
rect 2409 18819 2467 18825
rect 2409 18785 2421 18819
rect 2455 18785 2467 18819
rect 2409 18779 2467 18785
rect 2593 18819 2651 18825
rect 2593 18785 2605 18819
rect 2639 18816 2651 18819
rect 3326 18816 3332 18828
rect 2639 18788 2774 18816
rect 3287 18788 3332 18816
rect 2639 18785 2651 18788
rect 2593 18779 2651 18785
rect 2746 18612 2774 18788
rect 3326 18776 3332 18788
rect 3384 18776 3390 18828
rect 4908 18816 4936 18847
rect 5074 18844 5080 18856
rect 5132 18844 5138 18896
rect 8389 18887 8447 18893
rect 8389 18853 8401 18887
rect 8435 18884 8447 18887
rect 10962 18884 10968 18896
rect 8435 18856 10968 18884
rect 8435 18853 8447 18856
rect 8389 18847 8447 18853
rect 10962 18844 10968 18856
rect 11020 18844 11026 18896
rect 11256 18884 11284 18924
rect 11425 18921 11437 18955
rect 11471 18952 11483 18955
rect 11471 18924 16804 18952
rect 11471 18921 11483 18924
rect 11425 18915 11483 18921
rect 13449 18887 13507 18893
rect 13449 18884 13461 18887
rect 11256 18856 13461 18884
rect 13449 18853 13461 18856
rect 13495 18884 13507 18887
rect 15470 18884 15476 18896
rect 13495 18856 15476 18884
rect 13495 18853 13507 18856
rect 13449 18847 13507 18853
rect 15470 18844 15476 18856
rect 15528 18844 15534 18896
rect 16298 18884 16304 18896
rect 15764 18856 16304 18884
rect 5537 18819 5595 18825
rect 5537 18816 5549 18819
rect 4908 18788 5549 18816
rect 5537 18785 5549 18788
rect 5583 18785 5595 18819
rect 5537 18779 5595 18785
rect 5718 18776 5724 18828
rect 5776 18816 5782 18828
rect 6178 18816 6184 18828
rect 5776 18788 6184 18816
rect 5776 18776 5782 18788
rect 6178 18776 6184 18788
rect 6236 18776 6242 18828
rect 6822 18776 6828 18828
rect 6880 18816 6886 18828
rect 8297 18819 8355 18825
rect 8297 18816 8309 18819
rect 6880 18788 8309 18816
rect 6880 18776 6886 18788
rect 8297 18785 8309 18788
rect 8343 18785 8355 18819
rect 8478 18816 8484 18828
rect 8439 18788 8484 18816
rect 8297 18779 8355 18785
rect 8478 18776 8484 18788
rect 8536 18776 8542 18828
rect 9674 18816 9680 18828
rect 9635 18788 9680 18816
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 9861 18819 9919 18825
rect 9861 18785 9873 18819
rect 9907 18816 9919 18819
rect 10686 18816 10692 18828
rect 9907 18788 10692 18816
rect 9907 18785 9919 18788
rect 9861 18779 9919 18785
rect 10686 18776 10692 18788
rect 10744 18776 10750 18828
rect 10781 18819 10839 18825
rect 10781 18785 10793 18819
rect 10827 18816 10839 18819
rect 11330 18816 11336 18828
rect 10827 18788 11336 18816
rect 10827 18785 10839 18788
rect 10781 18779 10839 18785
rect 11330 18776 11336 18788
rect 11388 18776 11394 18828
rect 11514 18816 11520 18828
rect 11475 18788 11520 18816
rect 11514 18776 11520 18788
rect 11572 18776 11578 18828
rect 13354 18816 13360 18828
rect 12360 18788 13360 18816
rect 10226 18708 10232 18760
rect 10284 18748 10290 18760
rect 10505 18751 10563 18757
rect 10505 18748 10517 18751
rect 10284 18720 10517 18748
rect 10284 18708 10290 18720
rect 10505 18717 10517 18720
rect 10551 18717 10563 18751
rect 10505 18711 10563 18717
rect 10594 18708 10600 18760
rect 10652 18748 10658 18760
rect 11425 18751 11483 18757
rect 11425 18748 11437 18751
rect 10652 18720 11437 18748
rect 10652 18708 10658 18720
rect 11425 18717 11437 18720
rect 11471 18717 11483 18751
rect 11425 18711 11483 18717
rect 11698 18708 11704 18760
rect 11756 18748 11762 18760
rect 12360 18757 12388 18788
rect 13354 18776 13360 18788
rect 13412 18776 13418 18828
rect 13630 18816 13636 18828
rect 13591 18788 13636 18816
rect 13630 18776 13636 18788
rect 13688 18776 13694 18828
rect 13817 18819 13875 18825
rect 13817 18785 13829 18819
rect 13863 18816 13875 18819
rect 13906 18816 13912 18828
rect 13863 18788 13912 18816
rect 13863 18785 13875 18788
rect 13817 18779 13875 18785
rect 13906 18776 13912 18788
rect 13964 18816 13970 18828
rect 13964 18788 14320 18816
rect 13964 18776 13970 18788
rect 12345 18751 12403 18757
rect 12345 18748 12357 18751
rect 11756 18720 12357 18748
rect 11756 18708 11762 18720
rect 12345 18717 12357 18720
rect 12391 18717 12403 18751
rect 12345 18711 12403 18717
rect 12434 18708 12440 18760
rect 12492 18748 12498 18760
rect 12710 18748 12716 18760
rect 12492 18720 12537 18748
rect 12671 18720 12716 18748
rect 12492 18708 12498 18720
rect 12710 18708 12716 18720
rect 12768 18708 12774 18760
rect 12897 18751 12955 18757
rect 12897 18717 12909 18751
rect 12943 18748 12955 18751
rect 13538 18748 13544 18760
rect 12943 18720 13544 18748
rect 12943 18717 12955 18720
rect 12897 18711 12955 18717
rect 13538 18708 13544 18720
rect 13596 18708 13602 18760
rect 4062 18640 4068 18692
rect 4120 18680 4126 18692
rect 10318 18680 10324 18692
rect 4120 18652 10324 18680
rect 4120 18640 4126 18652
rect 10318 18640 10324 18652
rect 10376 18640 10382 18692
rect 10410 18640 10416 18692
rect 10468 18680 10474 18692
rect 14292 18680 14320 18788
rect 14918 18776 14924 18828
rect 14976 18816 14982 18828
rect 15764 18825 15792 18856
rect 16298 18844 16304 18856
rect 16356 18844 16362 18896
rect 16776 18893 16804 18924
rect 17402 18912 17408 18964
rect 17460 18952 17466 18964
rect 17770 18952 17776 18964
rect 17460 18924 17776 18952
rect 17460 18912 17466 18924
rect 17770 18912 17776 18924
rect 17828 18952 17834 18964
rect 17828 18924 19288 18952
rect 17828 18912 17834 18924
rect 16763 18887 16821 18893
rect 16763 18853 16775 18887
rect 16809 18853 16821 18887
rect 16763 18847 16821 18853
rect 18046 18844 18052 18896
rect 18104 18884 18110 18896
rect 19260 18884 19288 18924
rect 19886 18912 19892 18964
rect 19944 18952 19950 18964
rect 25130 18952 25136 18964
rect 19944 18924 25136 18952
rect 19944 18912 19950 18924
rect 25130 18912 25136 18924
rect 25188 18912 25194 18964
rect 26510 18952 26516 18964
rect 26068 18924 26516 18952
rect 26068 18884 26096 18924
rect 26510 18912 26516 18924
rect 26568 18912 26574 18964
rect 32122 18912 32128 18964
rect 32180 18952 32186 18964
rect 32677 18955 32735 18961
rect 32677 18952 32689 18955
rect 32180 18924 32689 18952
rect 32180 18912 32186 18924
rect 32677 18921 32689 18924
rect 32723 18921 32735 18955
rect 32677 18915 32735 18921
rect 33045 18955 33103 18961
rect 33045 18921 33057 18955
rect 33091 18952 33103 18955
rect 33594 18952 33600 18964
rect 33091 18924 33600 18952
rect 33091 18921 33103 18924
rect 33045 18915 33103 18921
rect 33594 18912 33600 18924
rect 33652 18912 33658 18964
rect 18104 18856 19196 18884
rect 19260 18856 20116 18884
rect 18104 18844 18110 18856
rect 15013 18819 15071 18825
rect 15013 18816 15025 18819
rect 14976 18788 15025 18816
rect 14976 18776 14982 18788
rect 15013 18785 15025 18788
rect 15059 18785 15071 18819
rect 15013 18779 15071 18785
rect 15749 18819 15807 18825
rect 15749 18785 15761 18819
rect 15795 18785 15807 18819
rect 15749 18779 15807 18785
rect 15933 18819 15991 18825
rect 15933 18785 15945 18819
rect 15979 18785 15991 18819
rect 15933 18779 15991 18785
rect 15194 18748 15200 18760
rect 15155 18720 15200 18748
rect 15194 18708 15200 18720
rect 15252 18708 15258 18760
rect 15948 18748 15976 18779
rect 16022 18776 16028 18828
rect 16080 18816 16086 18828
rect 19168 18825 19196 18856
rect 18785 18819 18843 18825
rect 18785 18816 18797 18819
rect 16080 18788 18797 18816
rect 16080 18776 16086 18788
rect 18785 18785 18797 18788
rect 18831 18785 18843 18819
rect 18785 18779 18843 18785
rect 19153 18819 19211 18825
rect 19153 18785 19165 18819
rect 19199 18816 19211 18819
rect 19702 18816 19708 18828
rect 19199 18788 19708 18816
rect 19199 18785 19211 18788
rect 19153 18779 19211 18785
rect 19702 18776 19708 18788
rect 19760 18776 19766 18828
rect 19886 18816 19892 18828
rect 19847 18788 19892 18816
rect 19886 18776 19892 18788
rect 19944 18776 19950 18828
rect 20088 18825 20116 18856
rect 25976 18856 26096 18884
rect 20073 18819 20131 18825
rect 20073 18785 20085 18819
rect 20119 18785 20131 18819
rect 20073 18779 20131 18785
rect 20162 18776 20168 18828
rect 20220 18816 20226 18828
rect 25225 18819 25283 18825
rect 20220 18788 20265 18816
rect 20220 18776 20226 18788
rect 25225 18785 25237 18819
rect 25271 18816 25283 18819
rect 25314 18816 25320 18828
rect 25271 18788 25320 18816
rect 25271 18785 25283 18788
rect 25225 18779 25283 18785
rect 25314 18776 25320 18788
rect 25372 18776 25378 18828
rect 25976 18825 26004 18856
rect 26326 18844 26332 18896
rect 26384 18884 26390 18896
rect 26789 18887 26847 18893
rect 26789 18884 26801 18887
rect 26384 18856 26801 18884
rect 26384 18844 26390 18856
rect 26789 18853 26801 18856
rect 26835 18884 26847 18887
rect 28721 18887 28779 18893
rect 28721 18884 28733 18887
rect 26835 18856 28733 18884
rect 26835 18853 26847 18856
rect 26789 18847 26847 18853
rect 28721 18853 28733 18856
rect 28767 18853 28779 18887
rect 30742 18884 30748 18896
rect 30703 18856 30748 18884
rect 28721 18847 28779 18853
rect 30742 18844 30748 18856
rect 30800 18844 30806 18896
rect 32582 18884 32588 18896
rect 31970 18856 32588 18884
rect 32582 18844 32588 18856
rect 32640 18844 32646 18896
rect 25961 18819 26019 18825
rect 25961 18785 25973 18819
rect 26007 18785 26019 18819
rect 26142 18816 26148 18828
rect 26103 18788 26148 18816
rect 25961 18779 26019 18785
rect 26142 18776 26148 18788
rect 26200 18776 26206 18828
rect 26694 18816 26700 18828
rect 26655 18788 26700 18816
rect 26694 18776 26700 18788
rect 26752 18776 26758 18828
rect 26973 18819 27031 18825
rect 26973 18785 26985 18819
rect 27019 18816 27031 18819
rect 27246 18816 27252 18828
rect 27019 18788 27252 18816
rect 27019 18785 27031 18788
rect 26973 18779 27031 18785
rect 27246 18776 27252 18788
rect 27304 18776 27310 18828
rect 28166 18816 28172 18828
rect 28127 18788 28172 18816
rect 28166 18776 28172 18788
rect 28224 18776 28230 18828
rect 28353 18819 28411 18825
rect 28353 18785 28365 18819
rect 28399 18816 28411 18819
rect 28442 18816 28448 18828
rect 28399 18788 28448 18816
rect 28399 18785 28411 18788
rect 28353 18779 28411 18785
rect 18966 18748 18972 18760
rect 15948 18720 17908 18748
rect 18927 18720 18972 18748
rect 17880 18692 17908 18720
rect 18966 18708 18972 18720
rect 19024 18708 19030 18760
rect 19610 18748 19616 18760
rect 19571 18720 19616 18748
rect 19610 18708 19616 18720
rect 19668 18708 19674 18760
rect 19794 18748 19800 18760
rect 19755 18720 19800 18748
rect 19794 18708 19800 18720
rect 19852 18708 19858 18760
rect 20346 18748 20352 18760
rect 20307 18720 20352 18748
rect 20346 18708 20352 18720
rect 20404 18708 20410 18760
rect 25501 18751 25559 18757
rect 25501 18717 25513 18751
rect 25547 18748 25559 18751
rect 26053 18751 26111 18757
rect 26053 18748 26065 18751
rect 25547 18720 26065 18748
rect 25547 18717 25559 18720
rect 25501 18711 25559 18717
rect 26053 18717 26065 18720
rect 26099 18717 26111 18751
rect 26712 18748 26740 18776
rect 28368 18748 28396 18779
rect 28442 18776 28448 18788
rect 28500 18776 28506 18828
rect 29822 18776 29828 18828
rect 29880 18816 29886 18828
rect 30469 18819 30527 18825
rect 30469 18816 30481 18819
rect 29880 18788 30481 18816
rect 29880 18776 29886 18788
rect 30469 18785 30481 18788
rect 30515 18785 30527 18819
rect 30469 18779 30527 18785
rect 26712 18720 28396 18748
rect 26053 18711 26111 18717
rect 31202 18708 31208 18760
rect 31260 18748 31266 18760
rect 32214 18748 32220 18760
rect 31260 18720 31800 18748
rect 32175 18720 32220 18748
rect 31260 18708 31266 18720
rect 16850 18680 16856 18692
rect 10468 18652 10548 18680
rect 14292 18652 16856 18680
rect 10468 18640 10474 18652
rect 3145 18615 3203 18621
rect 3145 18612 3157 18615
rect 2746 18584 3157 18612
rect 3145 18581 3157 18584
rect 3191 18612 3203 18615
rect 4893 18615 4951 18621
rect 4893 18612 4905 18615
rect 3191 18584 4905 18612
rect 3191 18581 3203 18584
rect 3145 18575 3203 18581
rect 4893 18581 4905 18584
rect 4939 18612 4951 18615
rect 5718 18612 5724 18624
rect 4939 18584 5724 18612
rect 4939 18581 4951 18584
rect 4893 18575 4951 18581
rect 5718 18572 5724 18584
rect 5776 18572 5782 18624
rect 10520 18612 10548 18652
rect 16850 18640 16856 18652
rect 16908 18640 16914 18692
rect 17862 18640 17868 18692
rect 17920 18680 17926 18692
rect 18785 18683 18843 18689
rect 18785 18680 18797 18683
rect 17920 18652 18797 18680
rect 17920 18640 17926 18652
rect 18785 18649 18797 18652
rect 18831 18649 18843 18683
rect 19518 18680 19524 18692
rect 18785 18643 18843 18649
rect 18984 18652 19524 18680
rect 10597 18615 10655 18621
rect 10597 18612 10609 18615
rect 10520 18584 10609 18612
rect 10597 18581 10609 18584
rect 10643 18581 10655 18615
rect 10597 18575 10655 18581
rect 10686 18572 10692 18624
rect 10744 18612 10750 18624
rect 11609 18615 11667 18621
rect 10744 18584 10789 18612
rect 10744 18572 10750 18584
rect 11609 18581 11621 18615
rect 11655 18612 11667 18615
rect 12802 18612 12808 18624
rect 11655 18584 12808 18612
rect 11655 18581 11667 18584
rect 11609 18575 11667 18581
rect 12802 18572 12808 18584
rect 12860 18572 12866 18624
rect 17034 18572 17040 18624
rect 17092 18612 17098 18624
rect 18049 18615 18107 18621
rect 18049 18612 18061 18615
rect 17092 18584 18061 18612
rect 17092 18572 17098 18584
rect 18049 18581 18061 18584
rect 18095 18612 18107 18615
rect 18984 18612 19012 18652
rect 19518 18640 19524 18652
rect 19576 18640 19582 18692
rect 25317 18683 25375 18689
rect 25317 18649 25329 18683
rect 25363 18680 25375 18683
rect 25958 18680 25964 18692
rect 25363 18652 25964 18680
rect 25363 18649 25375 18652
rect 25317 18643 25375 18649
rect 25958 18640 25964 18652
rect 26016 18640 26022 18692
rect 27890 18680 27896 18692
rect 27851 18652 27896 18680
rect 27890 18640 27896 18652
rect 27948 18640 27954 18692
rect 31772 18680 31800 18720
rect 32214 18708 32220 18720
rect 32272 18748 32278 18760
rect 33137 18751 33195 18757
rect 33137 18748 33149 18751
rect 32272 18720 33149 18748
rect 32272 18708 32278 18720
rect 33137 18717 33149 18720
rect 33183 18717 33195 18751
rect 33137 18711 33195 18717
rect 33229 18751 33287 18757
rect 33229 18717 33241 18751
rect 33275 18717 33287 18751
rect 33229 18711 33287 18717
rect 33244 18680 33272 18711
rect 31772 18652 33272 18680
rect 18095 18584 19012 18612
rect 18095 18581 18107 18584
rect 18049 18575 18107 18581
rect 19058 18572 19064 18624
rect 19116 18612 19122 18624
rect 19705 18615 19763 18621
rect 19705 18612 19717 18615
rect 19116 18584 19717 18612
rect 19116 18572 19122 18584
rect 19705 18581 19717 18584
rect 19751 18581 19763 18615
rect 19705 18575 19763 18581
rect 25406 18572 25412 18624
rect 25464 18612 25470 18624
rect 27154 18612 27160 18624
rect 25464 18584 25509 18612
rect 27115 18584 27160 18612
rect 25464 18572 25470 18584
rect 27154 18572 27160 18584
rect 27212 18572 27218 18624
rect 27985 18615 28043 18621
rect 27985 18581 27997 18615
rect 28031 18612 28043 18615
rect 28074 18612 28080 18624
rect 28031 18584 28080 18612
rect 28031 18581 28043 18584
rect 27985 18575 28043 18581
rect 28074 18572 28080 18584
rect 28132 18572 28138 18624
rect 1104 18522 34316 18544
rect 1104 18470 6517 18522
rect 6569 18470 6581 18522
rect 6633 18470 6645 18522
rect 6697 18470 6709 18522
rect 6761 18470 17588 18522
rect 17640 18470 17652 18522
rect 17704 18470 17716 18522
rect 17768 18470 17780 18522
rect 17832 18470 28658 18522
rect 28710 18470 28722 18522
rect 28774 18470 28786 18522
rect 28838 18470 28850 18522
rect 28902 18470 34316 18522
rect 1104 18448 34316 18470
rect 4065 18411 4123 18417
rect 4065 18377 4077 18411
rect 4111 18377 4123 18411
rect 4065 18371 4123 18377
rect 4080 18272 4108 18371
rect 8202 18368 8208 18420
rect 8260 18408 8266 18420
rect 9582 18408 9588 18420
rect 8260 18380 9588 18408
rect 8260 18368 8266 18380
rect 9582 18368 9588 18380
rect 9640 18368 9646 18420
rect 10686 18368 10692 18420
rect 10744 18408 10750 18420
rect 10873 18411 10931 18417
rect 10873 18408 10885 18411
rect 10744 18380 10885 18408
rect 10744 18368 10750 18380
rect 10873 18377 10885 18380
rect 10919 18377 10931 18411
rect 10873 18371 10931 18377
rect 10962 18368 10968 18420
rect 11020 18408 11026 18420
rect 12342 18408 12348 18420
rect 11020 18380 12348 18408
rect 11020 18368 11026 18380
rect 12342 18368 12348 18380
rect 12400 18368 12406 18420
rect 12434 18368 12440 18420
rect 12492 18408 12498 18420
rect 12894 18408 12900 18420
rect 12492 18380 12900 18408
rect 12492 18368 12498 18380
rect 12894 18368 12900 18380
rect 12952 18408 12958 18420
rect 15010 18408 15016 18420
rect 12952 18380 15016 18408
rect 12952 18368 12958 18380
rect 15010 18368 15016 18380
rect 15068 18368 15074 18420
rect 15746 18368 15752 18420
rect 15804 18408 15810 18420
rect 16301 18411 16359 18417
rect 16301 18408 16313 18411
rect 15804 18380 16313 18408
rect 15804 18368 15810 18380
rect 16301 18377 16313 18380
rect 16347 18377 16359 18411
rect 16301 18371 16359 18377
rect 17402 18368 17408 18420
rect 17460 18408 17466 18420
rect 17589 18411 17647 18417
rect 17589 18408 17601 18411
rect 17460 18380 17601 18408
rect 17460 18368 17466 18380
rect 17589 18377 17601 18380
rect 17635 18377 17647 18411
rect 19886 18408 19892 18420
rect 17589 18371 17647 18377
rect 17696 18380 19892 18408
rect 12250 18340 12256 18352
rect 9232 18312 12256 18340
rect 5074 18272 5080 18284
rect 4080 18244 5080 18272
rect 2498 18204 2504 18216
rect 2459 18176 2504 18204
rect 2498 18164 2504 18176
rect 2556 18164 2562 18216
rect 2685 18207 2743 18213
rect 2685 18173 2697 18207
rect 2731 18204 2743 18207
rect 2774 18204 2780 18216
rect 2731 18176 2780 18204
rect 2731 18173 2743 18176
rect 2685 18167 2743 18173
rect 2774 18164 2780 18176
rect 2832 18164 2838 18216
rect 2961 18207 3019 18213
rect 2961 18173 2973 18207
rect 3007 18204 3019 18207
rect 3234 18204 3240 18216
rect 3007 18176 3240 18204
rect 3007 18173 3019 18176
rect 2961 18167 3019 18173
rect 3234 18164 3240 18176
rect 3292 18164 3298 18216
rect 5000 18213 5028 18244
rect 5074 18232 5080 18244
rect 5132 18232 5138 18284
rect 5184 18244 6868 18272
rect 5184 18213 5212 18244
rect 6840 18216 6868 18244
rect 4893 18207 4951 18213
rect 4893 18204 4905 18207
rect 4172 18176 4905 18204
rect 3050 18136 3056 18148
rect 3011 18108 3056 18136
rect 3050 18096 3056 18108
rect 3108 18096 3114 18148
rect 4044 18139 4102 18145
rect 4044 18105 4056 18139
rect 4090 18136 4102 18139
rect 4172 18136 4200 18176
rect 4893 18173 4905 18176
rect 4939 18173 4951 18207
rect 4893 18167 4951 18173
rect 4985 18207 5043 18213
rect 4985 18173 4997 18207
rect 5031 18173 5043 18207
rect 4985 18167 5043 18173
rect 5169 18207 5227 18213
rect 5169 18173 5181 18207
rect 5215 18173 5227 18207
rect 5169 18167 5227 18173
rect 4090 18108 4200 18136
rect 4090 18105 4102 18108
rect 4044 18099 4102 18105
rect 4246 18096 4252 18148
rect 4304 18136 4310 18148
rect 4908 18136 4936 18167
rect 5258 18164 5264 18216
rect 5316 18204 5322 18216
rect 5316 18176 5361 18204
rect 5316 18164 5322 18176
rect 6822 18164 6828 18216
rect 6880 18204 6886 18216
rect 7101 18207 7159 18213
rect 7101 18204 7113 18207
rect 6880 18176 7113 18204
rect 6880 18164 6886 18176
rect 7101 18173 7113 18176
rect 7147 18173 7159 18207
rect 7101 18167 7159 18173
rect 7282 18164 7288 18216
rect 7340 18204 7346 18216
rect 9232 18213 9260 18312
rect 12250 18300 12256 18312
rect 12308 18300 12314 18352
rect 9858 18272 9864 18284
rect 9462 18244 9864 18272
rect 9462 18213 9490 18244
rect 9858 18232 9864 18244
rect 9916 18232 9922 18284
rect 12710 18272 12716 18284
rect 11072 18244 12296 18272
rect 7653 18207 7711 18213
rect 7653 18204 7665 18207
rect 7340 18176 7665 18204
rect 7340 18164 7346 18176
rect 7653 18173 7665 18176
rect 7699 18173 7711 18207
rect 7653 18167 7711 18173
rect 9125 18207 9183 18213
rect 9125 18173 9137 18207
rect 9171 18173 9183 18207
rect 9125 18167 9183 18173
rect 9217 18207 9275 18213
rect 9217 18173 9229 18207
rect 9263 18173 9275 18207
rect 9217 18167 9275 18173
rect 9427 18207 9490 18213
rect 9427 18173 9439 18207
rect 9473 18176 9490 18207
rect 9473 18173 9485 18176
rect 9427 18167 9485 18173
rect 6178 18136 6184 18148
rect 4304 18108 4349 18136
rect 4908 18108 6184 18136
rect 4304 18096 4310 18108
rect 6178 18096 6184 18108
rect 6236 18096 6242 18148
rect 6917 18139 6975 18145
rect 6917 18105 6929 18139
rect 6963 18105 6975 18139
rect 6917 18099 6975 18105
rect 3878 18068 3884 18080
rect 3839 18040 3884 18068
rect 3878 18028 3884 18040
rect 3936 18028 3942 18080
rect 4154 18028 4160 18080
rect 4212 18068 4218 18080
rect 4709 18071 4767 18077
rect 4709 18068 4721 18071
rect 4212 18040 4721 18068
rect 4212 18028 4218 18040
rect 4709 18037 4721 18040
rect 4755 18037 4767 18071
rect 4709 18031 4767 18037
rect 4982 18028 4988 18080
rect 5040 18068 5046 18080
rect 6932 18068 6960 18099
rect 5040 18040 6960 18068
rect 5040 18028 5046 18040
rect 8478 18028 8484 18080
rect 8536 18068 8542 18080
rect 8941 18071 8999 18077
rect 8941 18068 8953 18071
rect 8536 18040 8953 18068
rect 8536 18028 8542 18040
rect 8941 18037 8953 18040
rect 8987 18037 8999 18071
rect 9140 18068 9168 18167
rect 9582 18164 9588 18216
rect 9640 18204 9646 18216
rect 10229 18207 10287 18213
rect 9640 18176 9685 18204
rect 9640 18164 9646 18176
rect 10229 18173 10241 18207
rect 10275 18173 10287 18207
rect 10229 18167 10287 18173
rect 10321 18207 10379 18213
rect 10321 18173 10333 18207
rect 10367 18204 10379 18207
rect 11072 18204 11100 18244
rect 10367 18176 11100 18204
rect 10367 18173 10379 18176
rect 10321 18167 10379 18173
rect 9309 18139 9367 18145
rect 9309 18105 9321 18139
rect 9355 18136 9367 18139
rect 10042 18136 10048 18148
rect 9355 18108 10048 18136
rect 9355 18105 9367 18108
rect 9309 18099 9367 18105
rect 10042 18096 10048 18108
rect 10100 18096 10106 18148
rect 9950 18068 9956 18080
rect 9140 18040 9956 18068
rect 8941 18031 8999 18037
rect 9950 18028 9956 18040
rect 10008 18068 10014 18080
rect 10244 18068 10272 18167
rect 11146 18164 11152 18216
rect 11204 18204 11210 18216
rect 11204 18176 11249 18204
rect 11204 18164 11210 18176
rect 10873 18139 10931 18145
rect 10873 18105 10885 18139
rect 10919 18136 10931 18139
rect 12069 18139 12127 18145
rect 12069 18136 12081 18139
rect 10919 18108 12081 18136
rect 10919 18105 10931 18108
rect 10873 18099 10931 18105
rect 12069 18105 12081 18108
rect 12115 18105 12127 18139
rect 12069 18099 12127 18105
rect 11054 18068 11060 18080
rect 10008 18040 10272 18068
rect 11015 18040 11060 18068
rect 10008 18028 10014 18040
rect 11054 18028 11060 18040
rect 11112 18028 11118 18080
rect 12268 18068 12296 18244
rect 12360 18244 12716 18272
rect 12360 18213 12388 18244
rect 12710 18232 12716 18244
rect 12768 18232 12774 18284
rect 14826 18272 14832 18284
rect 14787 18244 14832 18272
rect 14826 18232 14832 18244
rect 14884 18232 14890 18284
rect 15764 18272 15792 18368
rect 16666 18300 16672 18352
rect 16724 18340 16730 18352
rect 17696 18340 17724 18380
rect 19886 18368 19892 18380
rect 19944 18368 19950 18420
rect 22646 18408 22652 18420
rect 20180 18380 22652 18408
rect 16724 18312 17724 18340
rect 16724 18300 16730 18312
rect 19702 18300 19708 18352
rect 19760 18340 19766 18352
rect 20180 18340 20208 18380
rect 22646 18368 22652 18380
rect 22704 18368 22710 18420
rect 26142 18368 26148 18420
rect 26200 18408 26206 18420
rect 26237 18411 26295 18417
rect 26237 18408 26249 18411
rect 26200 18380 26249 18408
rect 26200 18368 26206 18380
rect 26237 18377 26249 18380
rect 26283 18377 26295 18411
rect 27798 18408 27804 18420
rect 27759 18380 27804 18408
rect 26237 18371 26295 18377
rect 27798 18368 27804 18380
rect 27856 18368 27862 18420
rect 30558 18408 30564 18420
rect 30519 18380 30564 18408
rect 30558 18368 30564 18380
rect 30616 18408 30622 18420
rect 31570 18408 31576 18420
rect 30616 18380 31576 18408
rect 30616 18368 30622 18380
rect 31570 18368 31576 18380
rect 31628 18368 31634 18420
rect 19760 18312 20208 18340
rect 19760 18300 19766 18312
rect 20254 18300 20260 18352
rect 20312 18300 20318 18352
rect 18046 18272 18052 18284
rect 15028 18244 15792 18272
rect 16408 18244 18052 18272
rect 15028 18216 15056 18244
rect 12345 18207 12403 18213
rect 12345 18173 12357 18207
rect 12391 18173 12403 18207
rect 12345 18167 12403 18173
rect 12434 18164 12440 18216
rect 12492 18204 12498 18216
rect 12802 18204 12808 18216
rect 12492 18176 12537 18204
rect 12763 18176 12808 18204
rect 12492 18164 12498 18176
rect 12802 18164 12808 18176
rect 12860 18164 12866 18216
rect 13262 18204 13268 18216
rect 13223 18176 13268 18204
rect 13262 18164 13268 18176
rect 13320 18164 13326 18216
rect 13722 18204 13728 18216
rect 13683 18176 13728 18204
rect 13722 18164 13728 18176
rect 13780 18164 13786 18216
rect 15010 18204 15016 18216
rect 14923 18176 15016 18204
rect 15010 18164 15016 18176
rect 15068 18164 15074 18216
rect 15381 18207 15439 18213
rect 15381 18173 15393 18207
rect 15427 18173 15439 18207
rect 15381 18167 15439 18173
rect 15396 18080 15424 18167
rect 15470 18164 15476 18216
rect 15528 18204 15534 18216
rect 16408 18213 16436 18244
rect 18046 18232 18052 18244
rect 18104 18232 18110 18284
rect 19058 18272 19064 18284
rect 19019 18244 19064 18272
rect 19058 18232 19064 18244
rect 19116 18232 19122 18284
rect 19337 18275 19395 18281
rect 19337 18241 19349 18275
rect 19383 18272 19395 18275
rect 20272 18272 20300 18300
rect 21637 18275 21695 18281
rect 21637 18272 21649 18275
rect 19383 18244 21649 18272
rect 19383 18241 19395 18244
rect 19337 18235 19395 18241
rect 21637 18241 21649 18244
rect 21683 18272 21695 18275
rect 22738 18272 22744 18284
rect 21683 18244 22744 18272
rect 21683 18241 21695 18244
rect 21637 18235 21695 18241
rect 22738 18232 22744 18244
rect 22796 18232 22802 18284
rect 24397 18275 24455 18281
rect 24397 18241 24409 18275
rect 24443 18272 24455 18275
rect 24857 18275 24915 18281
rect 24857 18272 24869 18275
rect 24443 18244 24869 18272
rect 24443 18241 24455 18244
rect 24397 18235 24455 18241
rect 24857 18241 24869 18244
rect 24903 18241 24915 18275
rect 24857 18235 24915 18241
rect 16393 18207 16451 18213
rect 16393 18204 16405 18207
rect 15528 18176 16405 18204
rect 15528 18164 15534 18176
rect 16393 18173 16405 18176
rect 16439 18173 16451 18207
rect 16393 18167 16451 18173
rect 18598 18096 18604 18148
rect 18656 18096 18662 18148
rect 21082 18136 21088 18148
rect 20930 18108 21088 18136
rect 21082 18096 21088 18108
rect 21140 18096 21146 18148
rect 21358 18136 21364 18148
rect 21319 18108 21364 18136
rect 21358 18096 21364 18108
rect 21416 18096 21422 18148
rect 23658 18096 23664 18148
rect 23716 18096 23722 18148
rect 24118 18136 24124 18148
rect 24079 18108 24124 18136
rect 24118 18096 24124 18108
rect 24176 18096 24182 18148
rect 24872 18136 24900 18235
rect 27154 18232 27160 18284
rect 27212 18272 27218 18284
rect 27212 18244 28672 18272
rect 27212 18232 27218 18244
rect 25124 18207 25182 18213
rect 25124 18173 25136 18207
rect 25170 18204 25182 18207
rect 25406 18204 25412 18216
rect 25170 18176 25412 18204
rect 25170 18173 25182 18176
rect 25124 18167 25182 18173
rect 25406 18164 25412 18176
rect 25464 18164 25470 18216
rect 27798 18164 27804 18216
rect 27856 18204 27862 18216
rect 27893 18207 27951 18213
rect 27893 18204 27905 18207
rect 27856 18176 27905 18204
rect 27856 18164 27862 18176
rect 27893 18173 27905 18176
rect 27939 18173 27951 18207
rect 28074 18204 28080 18216
rect 28035 18176 28080 18204
rect 27893 18167 27951 18173
rect 28074 18164 28080 18176
rect 28132 18164 28138 18216
rect 28644 18213 28672 18244
rect 28629 18207 28687 18213
rect 28629 18173 28641 18207
rect 28675 18173 28687 18207
rect 28629 18167 28687 18173
rect 30377 18207 30435 18213
rect 30377 18173 30389 18207
rect 30423 18204 30435 18207
rect 30650 18204 30656 18216
rect 30423 18176 30656 18204
rect 30423 18173 30435 18176
rect 30377 18167 30435 18173
rect 30650 18164 30656 18176
rect 30708 18204 30714 18216
rect 30926 18204 30932 18216
rect 30708 18176 30932 18204
rect 30708 18164 30714 18176
rect 30926 18164 30932 18176
rect 30984 18164 30990 18216
rect 29822 18136 29828 18148
rect 24872 18108 29828 18136
rect 29822 18096 29828 18108
rect 29880 18096 29886 18148
rect 12710 18068 12716 18080
rect 12268 18040 12716 18068
rect 12710 18028 12716 18040
rect 12768 18028 12774 18080
rect 15378 18068 15384 18080
rect 15291 18040 15384 18068
rect 15378 18028 15384 18040
rect 15436 18068 15442 18080
rect 15838 18068 15844 18080
rect 15436 18040 15844 18068
rect 15436 18028 15442 18040
rect 15838 18028 15844 18040
rect 15896 18068 15902 18080
rect 18966 18068 18972 18080
rect 15896 18040 18972 18068
rect 15896 18028 15902 18040
rect 18966 18028 18972 18040
rect 19024 18068 19030 18080
rect 19889 18071 19947 18077
rect 19889 18068 19901 18071
rect 19024 18040 19901 18068
rect 19024 18028 19030 18040
rect 19889 18037 19901 18040
rect 19935 18068 19947 18071
rect 21266 18068 21272 18080
rect 19935 18040 21272 18068
rect 19935 18037 19947 18040
rect 19889 18031 19947 18037
rect 21266 18028 21272 18040
rect 21324 18028 21330 18080
rect 1104 17978 34316 18000
rect 1104 17926 12052 17978
rect 12104 17926 12116 17978
rect 12168 17926 12180 17978
rect 12232 17926 12244 17978
rect 12296 17926 23123 17978
rect 23175 17926 23187 17978
rect 23239 17926 23251 17978
rect 23303 17926 23315 17978
rect 23367 17926 34316 17978
rect 1104 17904 34316 17926
rect 1857 17867 1915 17873
rect 1857 17833 1869 17867
rect 1903 17864 1915 17867
rect 2498 17864 2504 17876
rect 1903 17836 2504 17864
rect 1903 17833 1915 17836
rect 1857 17827 1915 17833
rect 2498 17824 2504 17836
rect 2556 17824 2562 17876
rect 2866 17824 2872 17876
rect 2924 17864 2930 17876
rect 2961 17867 3019 17873
rect 2961 17864 2973 17867
rect 2924 17836 2973 17864
rect 2924 17824 2930 17836
rect 2961 17833 2973 17836
rect 3007 17833 3019 17867
rect 2961 17827 3019 17833
rect 8386 17824 8392 17876
rect 8444 17864 8450 17876
rect 9674 17864 9680 17876
rect 8444 17836 9680 17864
rect 8444 17824 8450 17836
rect 9674 17824 9680 17836
rect 9732 17864 9738 17876
rect 9732 17836 10824 17864
rect 9732 17824 9738 17836
rect 3050 17796 3056 17808
rect 3011 17768 3056 17796
rect 3050 17756 3056 17768
rect 3108 17756 3114 17808
rect 4706 17796 4712 17808
rect 4540 17768 4712 17796
rect 1765 17731 1823 17737
rect 1765 17697 1777 17731
rect 1811 17697 1823 17731
rect 1765 17691 1823 17697
rect 1949 17731 2007 17737
rect 1949 17697 1961 17731
rect 1995 17728 2007 17731
rect 2590 17728 2596 17740
rect 1995 17700 2596 17728
rect 1995 17697 2007 17700
rect 1949 17691 2007 17697
rect 1780 17660 1808 17691
rect 2590 17688 2596 17700
rect 2648 17688 2654 17740
rect 4338 17728 4344 17740
rect 4299 17700 4344 17728
rect 4338 17688 4344 17700
rect 4396 17688 4402 17740
rect 4540 17737 4568 17768
rect 4706 17756 4712 17768
rect 4764 17796 4770 17808
rect 5258 17796 5264 17808
rect 4764 17768 5264 17796
rect 4764 17756 4770 17768
rect 5258 17756 5264 17768
rect 5316 17756 5322 17808
rect 10796 17782 10824 17836
rect 17218 17824 17224 17876
rect 17276 17864 17282 17876
rect 17865 17867 17923 17873
rect 17865 17864 17877 17867
rect 17276 17836 17877 17864
rect 17276 17824 17282 17836
rect 17865 17833 17877 17836
rect 17911 17833 17923 17867
rect 17865 17827 17923 17833
rect 20809 17867 20867 17873
rect 20809 17833 20821 17867
rect 20855 17864 20867 17867
rect 21358 17864 21364 17876
rect 20855 17836 21364 17864
rect 20855 17833 20867 17836
rect 20809 17827 20867 17833
rect 21358 17824 21364 17836
rect 21416 17824 21422 17876
rect 22189 17867 22247 17873
rect 22189 17833 22201 17867
rect 22235 17864 22247 17867
rect 24118 17864 24124 17876
rect 22235 17836 24124 17864
rect 22235 17833 22247 17836
rect 22189 17827 22247 17833
rect 24118 17824 24124 17836
rect 24176 17824 24182 17876
rect 26605 17867 26663 17873
rect 26605 17833 26617 17867
rect 26651 17864 26663 17867
rect 27890 17864 27896 17876
rect 26651 17836 27896 17864
rect 26651 17833 26663 17836
rect 26605 17827 26663 17833
rect 27890 17824 27896 17836
rect 27948 17824 27954 17876
rect 12897 17799 12955 17805
rect 12897 17765 12909 17799
rect 12943 17796 12955 17799
rect 14918 17796 14924 17808
rect 12943 17768 14924 17796
rect 12943 17765 12955 17768
rect 12897 17759 12955 17765
rect 14918 17756 14924 17768
rect 14976 17756 14982 17808
rect 15378 17796 15384 17808
rect 15028 17768 15384 17796
rect 4525 17731 4583 17737
rect 4525 17697 4537 17731
rect 4571 17697 4583 17731
rect 4525 17691 4583 17697
rect 4985 17731 5043 17737
rect 4985 17697 4997 17731
rect 5031 17697 5043 17731
rect 5445 17731 5503 17737
rect 5445 17728 5457 17731
rect 4985 17691 5043 17697
rect 5368 17700 5457 17728
rect 2866 17660 2872 17672
rect 1780 17632 2872 17660
rect 2866 17620 2872 17632
rect 2924 17620 2930 17672
rect 4433 17663 4491 17669
rect 4433 17629 4445 17663
rect 4479 17660 4491 17663
rect 5000 17660 5028 17691
rect 4479 17632 5028 17660
rect 4479 17629 4491 17632
rect 4433 17623 4491 17629
rect 2501 17527 2559 17533
rect 2501 17493 2513 17527
rect 2547 17524 2559 17527
rect 2590 17524 2596 17536
rect 2547 17496 2596 17524
rect 2547 17493 2559 17496
rect 2501 17487 2559 17493
rect 2590 17484 2596 17496
rect 2648 17524 2654 17536
rect 4890 17524 4896 17536
rect 2648 17496 4896 17524
rect 2648 17484 2654 17496
rect 4890 17484 4896 17496
rect 4948 17524 4954 17536
rect 5368 17524 5396 17700
rect 5445 17697 5457 17700
rect 5491 17697 5503 17731
rect 5902 17728 5908 17740
rect 5863 17700 5908 17728
rect 5445 17691 5503 17697
rect 5902 17688 5908 17700
rect 5960 17688 5966 17740
rect 6178 17728 6184 17740
rect 6139 17700 6184 17728
rect 6178 17688 6184 17700
rect 6236 17688 6242 17740
rect 6362 17728 6368 17740
rect 6323 17700 6368 17728
rect 6362 17688 6368 17700
rect 6420 17688 6426 17740
rect 7466 17728 7472 17740
rect 7427 17700 7472 17728
rect 7466 17688 7472 17700
rect 7524 17688 7530 17740
rect 10410 17728 10416 17740
rect 10371 17700 10416 17728
rect 10410 17688 10416 17700
rect 10468 17688 10474 17740
rect 11882 17688 11888 17740
rect 11940 17728 11946 17740
rect 12805 17731 12863 17737
rect 12805 17728 12817 17731
rect 11940 17700 12817 17728
rect 11940 17688 11946 17700
rect 12805 17697 12817 17700
rect 12851 17697 12863 17731
rect 12805 17691 12863 17697
rect 12986 17688 12992 17740
rect 13044 17728 13050 17740
rect 13044 17700 13089 17728
rect 13044 17688 13050 17700
rect 14642 17688 14648 17740
rect 14700 17728 14706 17740
rect 14737 17731 14795 17737
rect 14737 17728 14749 17731
rect 14700 17700 14749 17728
rect 14700 17688 14706 17700
rect 14737 17697 14749 17700
rect 14783 17697 14795 17731
rect 14737 17691 14795 17697
rect 14829 17731 14887 17737
rect 14829 17697 14841 17731
rect 14875 17728 14887 17731
rect 15028 17728 15056 17768
rect 15378 17756 15384 17768
rect 15436 17756 15442 17808
rect 15841 17799 15899 17805
rect 15841 17765 15853 17799
rect 15887 17796 15899 17799
rect 15930 17796 15936 17808
rect 15887 17768 15936 17796
rect 15887 17765 15899 17768
rect 15841 17759 15899 17765
rect 15930 17756 15936 17768
rect 15988 17756 15994 17808
rect 16114 17756 16120 17808
rect 16172 17796 16178 17808
rect 22094 17796 22100 17808
rect 16172 17768 16330 17796
rect 21468 17768 22100 17796
rect 16172 17756 16178 17768
rect 14875 17700 15056 17728
rect 15105 17731 15163 17737
rect 14875 17697 14887 17700
rect 14829 17691 14887 17697
rect 15105 17697 15117 17731
rect 15151 17728 15163 17731
rect 15470 17728 15476 17740
rect 15151 17700 15476 17728
rect 15151 17697 15163 17700
rect 15105 17691 15163 17697
rect 15470 17688 15476 17700
rect 15528 17688 15534 17740
rect 17402 17688 17408 17740
rect 17460 17728 17466 17740
rect 17773 17731 17831 17737
rect 17773 17728 17785 17731
rect 17460 17700 17785 17728
rect 17460 17688 17466 17700
rect 17773 17697 17785 17700
rect 17819 17697 17831 17731
rect 17773 17691 17831 17697
rect 20533 17731 20591 17737
rect 20533 17697 20545 17731
rect 20579 17728 20591 17731
rect 20714 17728 20720 17740
rect 20579 17700 20720 17728
rect 20579 17697 20591 17700
rect 20533 17691 20591 17697
rect 20714 17688 20720 17700
rect 20772 17688 20778 17740
rect 21266 17728 21272 17740
rect 21227 17700 21272 17728
rect 21266 17688 21272 17700
rect 21324 17688 21330 17740
rect 21468 17737 21496 17768
rect 22094 17756 22100 17768
rect 22152 17796 22158 17808
rect 26786 17796 26792 17808
rect 22152 17768 22876 17796
rect 22152 17756 22158 17768
rect 22848 17740 22876 17768
rect 26528 17768 26792 17796
rect 21453 17731 21511 17737
rect 21453 17697 21465 17731
rect 21499 17697 21511 17731
rect 21453 17691 21511 17697
rect 21913 17731 21971 17737
rect 21913 17697 21925 17731
rect 21959 17697 21971 17731
rect 22646 17728 22652 17740
rect 22607 17700 22652 17728
rect 21913 17691 21971 17697
rect 10045 17663 10103 17669
rect 10045 17629 10057 17663
rect 10091 17660 10103 17663
rect 10778 17660 10784 17672
rect 10091 17632 10784 17660
rect 10091 17629 10103 17632
rect 10045 17623 10103 17629
rect 10778 17620 10784 17632
rect 10836 17620 10842 17672
rect 12529 17663 12587 17669
rect 12529 17629 12541 17663
rect 12575 17629 12587 17663
rect 12529 17623 12587 17629
rect 12621 17663 12679 17669
rect 12621 17629 12633 17663
rect 12667 17660 12679 17663
rect 12710 17660 12716 17672
rect 12667 17632 12716 17660
rect 12667 17629 12679 17632
rect 12621 17623 12679 17629
rect 6457 17595 6515 17601
rect 6457 17561 6469 17595
rect 6503 17592 6515 17595
rect 7190 17592 7196 17604
rect 6503 17564 7196 17592
rect 6503 17561 6515 17564
rect 6457 17555 6515 17561
rect 7190 17552 7196 17564
rect 7248 17552 7254 17604
rect 11606 17552 11612 17604
rect 11664 17592 11670 17604
rect 12544 17592 12572 17623
rect 12710 17620 12716 17632
rect 12768 17660 12774 17672
rect 13722 17660 13728 17672
rect 12768 17632 13728 17660
rect 12768 17620 12774 17632
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 15194 17620 15200 17672
rect 15252 17660 15258 17672
rect 15565 17663 15623 17669
rect 15565 17660 15577 17663
rect 15252 17632 15577 17660
rect 15252 17620 15258 17632
rect 15565 17629 15577 17632
rect 15611 17629 15623 17663
rect 17420 17660 17448 17688
rect 15565 17623 15623 17629
rect 15672 17632 17448 17660
rect 20809 17663 20867 17669
rect 15672 17592 15700 17632
rect 20809 17629 20821 17663
rect 20855 17660 20867 17663
rect 21361 17663 21419 17669
rect 21361 17660 21373 17663
rect 20855 17632 21373 17660
rect 20855 17629 20867 17632
rect 20809 17623 20867 17629
rect 21361 17629 21373 17632
rect 21407 17629 21419 17663
rect 21361 17623 21419 17629
rect 11664 17564 15700 17592
rect 21928 17592 21956 17691
rect 22646 17688 22652 17700
rect 22704 17688 22710 17740
rect 22830 17728 22836 17740
rect 22791 17700 22836 17728
rect 22830 17688 22836 17700
rect 22888 17688 22894 17740
rect 26528 17737 26556 17768
rect 26786 17756 26792 17768
rect 26844 17756 26850 17808
rect 27614 17796 27620 17808
rect 27356 17768 27620 17796
rect 27356 17737 27384 17768
rect 27614 17756 27620 17768
rect 27672 17756 27678 17808
rect 32582 17756 32588 17808
rect 32640 17756 32646 17808
rect 26513 17731 26571 17737
rect 26513 17697 26525 17731
rect 26559 17697 26571 17731
rect 26513 17691 26571 17697
rect 26697 17731 26755 17737
rect 26697 17697 26709 17731
rect 26743 17728 26755 17731
rect 27341 17731 27399 17737
rect 27341 17728 27353 17731
rect 26743 17700 27353 17728
rect 26743 17697 26755 17700
rect 26697 17691 26755 17697
rect 27341 17697 27353 17700
rect 27387 17697 27399 17731
rect 27982 17728 27988 17740
rect 27943 17700 27988 17728
rect 27341 17691 27399 17697
rect 22189 17663 22247 17669
rect 22189 17629 22201 17663
rect 22235 17660 22247 17663
rect 22741 17663 22799 17669
rect 22741 17660 22753 17663
rect 22235 17632 22753 17660
rect 22235 17629 22247 17632
rect 22189 17623 22247 17629
rect 22741 17629 22753 17632
rect 22787 17629 22799 17663
rect 22741 17623 22799 17629
rect 26418 17620 26424 17672
rect 26476 17660 26482 17672
rect 26528 17660 26556 17691
rect 27982 17688 27988 17700
rect 28040 17688 28046 17740
rect 31754 17688 31760 17740
rect 31812 17728 31818 17740
rect 31849 17731 31907 17737
rect 31849 17728 31861 17731
rect 31812 17700 31861 17728
rect 31812 17688 31818 17700
rect 31849 17697 31861 17700
rect 31895 17697 31907 17731
rect 31849 17691 31907 17697
rect 27249 17663 27307 17669
rect 27249 17660 27261 17663
rect 26476 17632 27261 17660
rect 26476 17620 26482 17632
rect 27249 17629 27261 17632
rect 27295 17629 27307 17663
rect 27798 17660 27804 17672
rect 27759 17632 27804 17660
rect 27249 17623 27307 17629
rect 27798 17620 27804 17632
rect 27856 17620 27862 17672
rect 28258 17660 28264 17672
rect 28219 17632 28264 17660
rect 28258 17620 28264 17632
rect 28316 17620 28322 17672
rect 32122 17660 32128 17672
rect 32083 17632 32128 17660
rect 32122 17620 32128 17632
rect 32180 17620 32186 17672
rect 21928 17564 22784 17592
rect 11664 17552 11670 17564
rect 22756 17536 22784 17564
rect 7374 17524 7380 17536
rect 4948 17496 5396 17524
rect 7335 17496 7380 17524
rect 4948 17484 4954 17496
rect 7374 17484 7380 17496
rect 7432 17484 7438 17536
rect 9582 17484 9588 17536
rect 9640 17524 9646 17536
rect 11514 17524 11520 17536
rect 9640 17496 11520 17524
rect 9640 17484 9646 17496
rect 11514 17484 11520 17496
rect 11572 17484 11578 17536
rect 11790 17524 11796 17536
rect 11749 17496 11796 17524
rect 11790 17484 11796 17496
rect 11848 17533 11854 17536
rect 11848 17527 11897 17533
rect 11848 17493 11851 17527
rect 11885 17524 11897 17527
rect 12342 17524 12348 17536
rect 11885 17496 12348 17524
rect 11885 17493 11897 17496
rect 11848 17487 11897 17493
rect 11848 17484 11854 17487
rect 12342 17484 12348 17496
rect 12400 17484 12406 17536
rect 13078 17484 13084 17536
rect 13136 17524 13142 17536
rect 13265 17527 13323 17533
rect 13265 17524 13277 17527
rect 13136 17496 13277 17524
rect 13136 17484 13142 17496
rect 13265 17493 13277 17496
rect 13311 17493 13323 17527
rect 13265 17487 13323 17493
rect 13630 17484 13636 17536
rect 13688 17524 13694 17536
rect 14826 17524 14832 17536
rect 13688 17496 14832 17524
rect 13688 17484 13694 17496
rect 14826 17484 14832 17496
rect 14884 17484 14890 17536
rect 17218 17484 17224 17536
rect 17276 17524 17282 17536
rect 17313 17527 17371 17533
rect 17313 17524 17325 17527
rect 17276 17496 17325 17524
rect 17276 17484 17282 17496
rect 17313 17493 17325 17496
rect 17359 17493 17371 17527
rect 17313 17487 17371 17493
rect 19610 17484 19616 17536
rect 19668 17524 19674 17536
rect 19978 17524 19984 17536
rect 19668 17496 19984 17524
rect 19668 17484 19674 17496
rect 19978 17484 19984 17496
rect 20036 17524 20042 17536
rect 20625 17527 20683 17533
rect 20625 17524 20637 17527
rect 20036 17496 20637 17524
rect 20036 17484 20042 17496
rect 20625 17493 20637 17496
rect 20671 17524 20683 17527
rect 22005 17527 22063 17533
rect 22005 17524 22017 17527
rect 20671 17496 22017 17524
rect 20671 17493 20683 17496
rect 20625 17487 20683 17493
rect 22005 17493 22017 17496
rect 22051 17493 22063 17527
rect 22005 17487 22063 17493
rect 22738 17484 22744 17536
rect 22796 17484 22802 17536
rect 33502 17484 33508 17536
rect 33560 17524 33566 17536
rect 33597 17527 33655 17533
rect 33597 17524 33609 17527
rect 33560 17496 33609 17524
rect 33560 17484 33566 17496
rect 33597 17493 33609 17496
rect 33643 17493 33655 17527
rect 33597 17487 33655 17493
rect 1104 17434 34316 17456
rect 1104 17382 6517 17434
rect 6569 17382 6581 17434
rect 6633 17382 6645 17434
rect 6697 17382 6709 17434
rect 6761 17382 17588 17434
rect 17640 17382 17652 17434
rect 17704 17382 17716 17434
rect 17768 17382 17780 17434
rect 17832 17382 28658 17434
rect 28710 17382 28722 17434
rect 28774 17382 28786 17434
rect 28838 17382 28850 17434
rect 28902 17382 34316 17434
rect 1104 17360 34316 17382
rect 2774 17280 2780 17332
rect 2832 17320 2838 17332
rect 4706 17320 4712 17332
rect 2832 17292 2877 17320
rect 4667 17292 4712 17320
rect 2832 17280 2838 17292
rect 4706 17280 4712 17292
rect 4764 17280 4770 17332
rect 4890 17320 4896 17332
rect 4851 17292 4896 17320
rect 4890 17280 4896 17292
rect 4948 17280 4954 17332
rect 5721 17323 5779 17329
rect 5721 17289 5733 17323
rect 5767 17320 5779 17323
rect 5902 17320 5908 17332
rect 5767 17292 5908 17320
rect 5767 17289 5779 17292
rect 5721 17283 5779 17289
rect 5902 17280 5908 17292
rect 5960 17280 5966 17332
rect 9950 17320 9956 17332
rect 8128 17292 9536 17320
rect 9911 17292 9956 17320
rect 7374 17184 7380 17196
rect 7335 17156 7380 17184
rect 7374 17144 7380 17156
rect 7432 17144 7438 17196
rect 2501 17119 2559 17125
rect 2501 17085 2513 17119
rect 2547 17085 2559 17119
rect 2501 17079 2559 17085
rect 2516 17048 2544 17079
rect 2590 17076 2596 17128
rect 2648 17116 2654 17128
rect 2648 17088 2693 17116
rect 2648 17076 2654 17088
rect 4246 17076 4252 17128
rect 4304 17116 4310 17128
rect 4798 17116 4804 17128
rect 4304 17088 4804 17116
rect 4304 17076 4310 17088
rect 4798 17076 4804 17088
rect 4856 17116 4862 17128
rect 5169 17119 5227 17125
rect 5169 17116 5181 17119
rect 4856 17088 5181 17116
rect 4856 17076 4862 17088
rect 5169 17085 5181 17088
rect 5215 17085 5227 17119
rect 5626 17116 5632 17128
rect 5587 17088 5632 17116
rect 5169 17079 5227 17085
rect 2866 17048 2872 17060
rect 2516 17020 2872 17048
rect 2866 17008 2872 17020
rect 2924 17008 2930 17060
rect 5184 17048 5212 17079
rect 5626 17076 5632 17088
rect 5684 17076 5690 17128
rect 5813 17119 5871 17125
rect 5813 17085 5825 17119
rect 5859 17085 5871 17119
rect 7190 17116 7196 17128
rect 7103 17088 7196 17116
rect 5813 17079 5871 17085
rect 5828 17048 5856 17079
rect 7190 17076 7196 17088
rect 7248 17116 7254 17128
rect 8128 17116 8156 17292
rect 9508 17252 9536 17292
rect 9950 17280 9956 17292
rect 10008 17280 10014 17332
rect 11146 17320 11152 17332
rect 11107 17292 11152 17320
rect 11146 17280 11152 17292
rect 11204 17280 11210 17332
rect 25130 17320 25136 17332
rect 12406 17292 25136 17320
rect 12406 17252 12434 17292
rect 25130 17280 25136 17292
rect 25188 17280 25194 17332
rect 28077 17323 28135 17329
rect 28077 17289 28089 17323
rect 28123 17320 28135 17323
rect 28166 17320 28172 17332
rect 28123 17292 28172 17320
rect 28123 17289 28135 17292
rect 28077 17283 28135 17289
rect 28166 17280 28172 17292
rect 28224 17280 28230 17332
rect 9508 17224 12434 17252
rect 13722 17212 13728 17264
rect 13780 17252 13786 17264
rect 30282 17252 30288 17264
rect 13780 17224 15240 17252
rect 13780 17212 13786 17224
rect 8478 17184 8484 17196
rect 8439 17156 8484 17184
rect 8478 17144 8484 17156
rect 8536 17144 8542 17196
rect 10781 17187 10839 17193
rect 10781 17153 10793 17187
rect 10827 17184 10839 17187
rect 11698 17184 11704 17196
rect 10827 17156 11704 17184
rect 10827 17153 10839 17156
rect 10781 17147 10839 17153
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 14737 17187 14795 17193
rect 14737 17184 14749 17187
rect 13464 17156 14749 17184
rect 7248 17088 8156 17116
rect 8205 17119 8263 17125
rect 7248 17076 7254 17088
rect 8205 17085 8217 17119
rect 8251 17085 8263 17119
rect 8205 17079 8263 17085
rect 10965 17119 11023 17125
rect 10965 17085 10977 17119
rect 11011 17085 11023 17119
rect 12526 17116 12532 17128
rect 12487 17088 12532 17116
rect 10965 17079 11023 17085
rect 5184 17020 5856 17048
rect 6362 17008 6368 17060
rect 6420 17048 6426 17060
rect 8220 17048 8248 17079
rect 6420 17020 8248 17048
rect 6420 17008 6426 17020
rect 8386 17008 8392 17060
rect 8444 17048 8450 17060
rect 8444 17020 8970 17048
rect 8444 17008 8450 17020
rect 6822 16980 6828 16992
rect 6783 16952 6828 16980
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 7282 16940 7288 16992
rect 7340 16980 7346 16992
rect 10980 16980 11008 17079
rect 12526 17076 12532 17088
rect 12584 17076 12590 17128
rect 13078 17116 13084 17128
rect 13039 17088 13084 17116
rect 13078 17076 13084 17088
rect 13136 17076 13142 17128
rect 13464 17125 13492 17156
rect 14737 17153 14749 17156
rect 14783 17153 14795 17187
rect 15102 17184 15108 17196
rect 15063 17156 15108 17184
rect 14737 17147 14795 17153
rect 15102 17144 15108 17156
rect 15160 17144 15166 17196
rect 15212 17193 15240 17224
rect 25424 17224 26096 17252
rect 30195 17224 30288 17252
rect 15197 17187 15255 17193
rect 15197 17153 15209 17187
rect 15243 17153 15255 17187
rect 15197 17147 15255 17153
rect 16114 17144 16120 17196
rect 16172 17184 16178 17196
rect 17310 17184 17316 17196
rect 16172 17156 17316 17184
rect 16172 17144 16178 17156
rect 17310 17144 17316 17156
rect 17368 17144 17374 17196
rect 21637 17187 21695 17193
rect 21637 17184 21649 17187
rect 17512 17156 19748 17184
rect 13449 17119 13507 17125
rect 13449 17085 13461 17119
rect 13495 17085 13507 17119
rect 13630 17116 13636 17128
rect 13591 17088 13636 17116
rect 13449 17079 13507 17085
rect 13630 17076 13636 17088
rect 13688 17076 13694 17128
rect 14001 17119 14059 17125
rect 14001 17085 14013 17119
rect 14047 17085 14059 17119
rect 14001 17079 14059 17085
rect 14921 17119 14979 17125
rect 14921 17085 14933 17119
rect 14967 17085 14979 17119
rect 14921 17079 14979 17085
rect 12434 17008 12440 17060
rect 12492 17048 12498 17060
rect 12492 17020 12537 17048
rect 12492 17008 12498 17020
rect 13538 17008 13544 17060
rect 13596 17048 13602 17060
rect 14016 17048 14044 17079
rect 13596 17020 14044 17048
rect 14936 17048 14964 17079
rect 15010 17076 15016 17128
rect 15068 17116 15074 17128
rect 15068 17088 15113 17116
rect 15068 17076 15074 17088
rect 15378 17048 15384 17060
rect 14936 17020 15384 17048
rect 13596 17008 13602 17020
rect 15378 17008 15384 17020
rect 15436 17008 15442 17060
rect 15746 17048 15752 17060
rect 15707 17020 15752 17048
rect 15746 17008 15752 17020
rect 15804 17008 15810 17060
rect 16117 17051 16175 17057
rect 16117 17017 16129 17051
rect 16163 17048 16175 17051
rect 17218 17048 17224 17060
rect 16163 17020 17224 17048
rect 16163 17017 16175 17020
rect 16117 17011 16175 17017
rect 17218 17008 17224 17020
rect 17276 17008 17282 17060
rect 12802 16980 12808 16992
rect 7340 16952 7385 16980
rect 10980 16952 12808 16980
rect 7340 16940 7346 16952
rect 12802 16940 12808 16952
rect 12860 16980 12866 16992
rect 13446 16980 13452 16992
rect 12860 16952 13452 16980
rect 12860 16940 12866 16952
rect 13446 16940 13452 16952
rect 13504 16980 13510 16992
rect 15764 16980 15792 17008
rect 13504 16952 15792 16980
rect 13504 16940 13510 16952
rect 17126 16940 17132 16992
rect 17184 16980 17190 16992
rect 17512 16989 17540 17156
rect 19720 17125 19748 17156
rect 19996 17156 21649 17184
rect 19996 17128 20024 17156
rect 21637 17153 21649 17156
rect 21683 17153 21695 17187
rect 21637 17147 21695 17153
rect 24578 17144 24584 17196
rect 24636 17184 24642 17196
rect 25424 17184 25452 17224
rect 25590 17184 25596 17196
rect 24636 17156 25452 17184
rect 25551 17156 25596 17184
rect 24636 17144 24642 17156
rect 25590 17144 25596 17156
rect 25648 17144 25654 17196
rect 26068 17193 26096 17224
rect 26053 17187 26111 17193
rect 26053 17153 26065 17187
rect 26099 17153 26111 17187
rect 26053 17147 26111 17153
rect 19245 17119 19303 17125
rect 19245 17085 19257 17119
rect 19291 17085 19303 17119
rect 19245 17079 19303 17085
rect 19705 17119 19763 17125
rect 19705 17085 19717 17119
rect 19751 17085 19763 17119
rect 19705 17079 19763 17085
rect 19889 17119 19947 17125
rect 19889 17085 19901 17119
rect 19935 17116 19947 17119
rect 19978 17116 19984 17128
rect 19935 17088 19984 17116
rect 19935 17085 19947 17088
rect 19889 17079 19947 17085
rect 18966 17048 18972 17060
rect 17497 16983 17555 16989
rect 17497 16980 17509 16983
rect 17184 16952 17509 16980
rect 17184 16940 17190 16952
rect 17497 16949 17509 16952
rect 17543 16949 17555 16983
rect 18524 16980 18552 17034
rect 18927 17020 18972 17048
rect 18966 17008 18972 17020
rect 19024 17008 19030 17060
rect 19260 17048 19288 17079
rect 19978 17076 19984 17088
rect 20036 17076 20042 17128
rect 21453 17119 21511 17125
rect 21453 17085 21465 17119
rect 21499 17116 21511 17119
rect 22094 17116 22100 17128
rect 21499 17088 22100 17116
rect 21499 17085 21511 17088
rect 21453 17079 21511 17085
rect 22094 17076 22100 17088
rect 22152 17076 22158 17128
rect 24946 17076 24952 17128
rect 25004 17116 25010 17128
rect 25685 17119 25743 17125
rect 25004 17088 25049 17116
rect 25004 17076 25010 17088
rect 25685 17085 25697 17119
rect 25731 17116 25743 17119
rect 26234 17116 26240 17128
rect 25731 17088 26240 17116
rect 25731 17085 25743 17088
rect 25685 17079 25743 17085
rect 26234 17076 26240 17088
rect 26292 17076 26298 17128
rect 26513 17119 26571 17125
rect 26513 17085 26525 17119
rect 26559 17085 26571 17119
rect 26694 17116 26700 17128
rect 26655 17088 26700 17116
rect 26513 17079 26571 17085
rect 20898 17048 20904 17060
rect 19260 17020 20904 17048
rect 20898 17008 20904 17020
rect 20956 17008 20962 17060
rect 23658 17008 23664 17060
rect 23716 17008 23722 17060
rect 24673 17051 24731 17057
rect 24673 17017 24685 17051
rect 24719 17017 24731 17051
rect 25958 17048 25964 17060
rect 25919 17020 25964 17048
rect 24673 17011 24731 17017
rect 18598 16980 18604 16992
rect 18524 16952 18604 16980
rect 17497 16943 17555 16949
rect 18598 16940 18604 16952
rect 18656 16940 18662 16992
rect 19794 16980 19800 16992
rect 19755 16952 19800 16980
rect 19794 16940 19800 16952
rect 19852 16940 19858 16992
rect 23201 16983 23259 16989
rect 23201 16949 23213 16983
rect 23247 16980 23259 16983
rect 23750 16980 23756 16992
rect 23247 16952 23756 16980
rect 23247 16949 23259 16952
rect 23201 16943 23259 16949
rect 23750 16940 23756 16952
rect 23808 16980 23814 16992
rect 24578 16980 24584 16992
rect 23808 16952 24584 16980
rect 23808 16940 23814 16952
rect 24578 16940 24584 16952
rect 24636 16940 24642 16992
rect 24688 16980 24716 17011
rect 25958 17008 25964 17020
rect 26016 17008 26022 17060
rect 26528 17048 26556 17079
rect 26694 17076 26700 17088
rect 26752 17076 26758 17128
rect 27982 17116 27988 17128
rect 27943 17088 27988 17116
rect 27982 17076 27988 17088
rect 28040 17076 28046 17128
rect 28169 17119 28227 17125
rect 28169 17085 28181 17119
rect 28215 17116 28227 17119
rect 28258 17116 28264 17128
rect 28215 17088 28264 17116
rect 28215 17085 28227 17088
rect 28169 17079 28227 17085
rect 28258 17076 28264 17088
rect 28316 17076 28322 17128
rect 28813 17119 28871 17125
rect 28813 17085 28825 17119
rect 28859 17085 28871 17119
rect 30208 17102 30236 17224
rect 30282 17212 30288 17224
rect 30340 17252 30346 17264
rect 32582 17252 32588 17264
rect 30340 17224 32588 17252
rect 30340 17212 30346 17224
rect 32582 17212 32588 17224
rect 32640 17212 32646 17264
rect 30558 17184 30564 17196
rect 30471 17156 30564 17184
rect 30558 17144 30564 17156
rect 30616 17184 30622 17196
rect 31389 17187 31447 17193
rect 31389 17184 31401 17187
rect 30616 17156 31401 17184
rect 30616 17144 30622 17156
rect 31389 17153 31401 17156
rect 31435 17153 31447 17187
rect 31389 17147 31447 17153
rect 31202 17116 31208 17128
rect 31163 17088 31208 17116
rect 28813 17079 28871 17085
rect 26068 17020 26556 17048
rect 25409 16983 25467 16989
rect 25409 16980 25421 16983
rect 24688 16952 25421 16980
rect 25409 16949 25421 16952
rect 25455 16949 25467 16983
rect 25409 16943 25467 16949
rect 25682 16940 25688 16992
rect 25740 16980 25746 16992
rect 26068 16980 26096 17020
rect 25740 16952 26096 16980
rect 25740 16940 25746 16952
rect 26142 16940 26148 16992
rect 26200 16980 26206 16992
rect 26513 16983 26571 16989
rect 26513 16980 26525 16983
rect 26200 16952 26525 16980
rect 26200 16940 26206 16952
rect 26513 16949 26525 16952
rect 26559 16949 26571 16983
rect 28828 16980 28856 17079
rect 31202 17076 31208 17088
rect 31260 17076 31266 17128
rect 31849 17119 31907 17125
rect 31849 17085 31861 17119
rect 31895 17085 31907 17119
rect 32030 17116 32036 17128
rect 31991 17088 32036 17116
rect 31849 17079 31907 17085
rect 29086 17048 29092 17060
rect 29047 17020 29092 17048
rect 29086 17008 29092 17020
rect 29144 17008 29150 17060
rect 30834 17008 30840 17060
rect 30892 17048 30898 17060
rect 31864 17048 31892 17079
rect 32030 17076 32036 17088
rect 32088 17076 32094 17128
rect 33134 17076 33140 17128
rect 33192 17116 33198 17128
rect 33413 17119 33471 17125
rect 33413 17116 33425 17119
rect 33192 17088 33425 17116
rect 33192 17076 33198 17088
rect 33413 17085 33425 17088
rect 33459 17085 33471 17119
rect 33413 17079 33471 17085
rect 32214 17048 32220 17060
rect 30892 17020 32220 17048
rect 30892 17008 30898 17020
rect 32214 17008 32220 17020
rect 32272 17008 32278 17060
rect 33594 17048 33600 17060
rect 33555 17020 33600 17048
rect 33594 17008 33600 17020
rect 33652 17008 33658 17060
rect 28994 16980 29000 16992
rect 28828 16952 29000 16980
rect 26513 16943 26571 16949
rect 28994 16940 29000 16952
rect 29052 16940 29058 16992
rect 31018 16980 31024 16992
rect 30979 16952 31024 16980
rect 31018 16940 31024 16952
rect 31076 16940 31082 16992
rect 31938 16980 31944 16992
rect 31899 16952 31944 16980
rect 31938 16940 31944 16952
rect 31996 16940 32002 16992
rect 1104 16890 34316 16912
rect 1104 16838 12052 16890
rect 12104 16838 12116 16890
rect 12168 16838 12180 16890
rect 12232 16838 12244 16890
rect 12296 16838 23123 16890
rect 23175 16838 23187 16890
rect 23239 16838 23251 16890
rect 23303 16838 23315 16890
rect 23367 16838 34316 16890
rect 1104 16816 34316 16838
rect 4338 16736 4344 16788
rect 4396 16776 4402 16788
rect 5537 16779 5595 16785
rect 5537 16776 5549 16779
rect 4396 16748 5549 16776
rect 4396 16736 4402 16748
rect 5537 16745 5549 16748
rect 5583 16745 5595 16779
rect 5537 16739 5595 16745
rect 7282 16736 7288 16788
rect 7340 16776 7346 16788
rect 7929 16779 7987 16785
rect 7929 16776 7941 16779
rect 7340 16748 7941 16776
rect 7340 16736 7346 16748
rect 7929 16745 7941 16748
rect 7975 16745 7987 16779
rect 11882 16776 11888 16788
rect 11843 16748 11888 16776
rect 7929 16739 7987 16745
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 12526 16776 12532 16788
rect 12487 16748 12532 16776
rect 12526 16736 12532 16748
rect 12584 16736 12590 16788
rect 14829 16779 14887 16785
rect 14829 16745 14841 16779
rect 14875 16776 14887 16779
rect 15102 16776 15108 16788
rect 14875 16748 15108 16776
rect 14875 16745 14887 16748
rect 14829 16739 14887 16745
rect 15102 16736 15108 16748
rect 15160 16736 15166 16788
rect 15749 16779 15807 16785
rect 15749 16745 15761 16779
rect 15795 16745 15807 16779
rect 17402 16776 17408 16788
rect 15749 16739 15807 16745
rect 15856 16748 17408 16776
rect 3053 16711 3111 16717
rect 3053 16677 3065 16711
rect 3099 16708 3111 16711
rect 3418 16708 3424 16720
rect 3099 16680 3424 16708
rect 3099 16677 3111 16680
rect 3053 16671 3111 16677
rect 3418 16668 3424 16680
rect 3476 16668 3482 16720
rect 6822 16717 6828 16720
rect 6816 16708 6828 16717
rect 6783 16680 6828 16708
rect 6816 16671 6828 16680
rect 6822 16668 6828 16671
rect 6880 16668 6886 16720
rect 2958 16649 2964 16652
rect 2956 16603 2964 16649
rect 3016 16640 3022 16652
rect 3145 16643 3203 16649
rect 3016 16612 3056 16640
rect 2958 16600 2964 16603
rect 3016 16600 3022 16612
rect 3145 16609 3157 16643
rect 3191 16609 3203 16643
rect 3326 16640 3332 16652
rect 3287 16612 3332 16640
rect 3145 16603 3203 16609
rect 3160 16572 3188 16603
rect 3326 16600 3332 16612
rect 3384 16600 3390 16652
rect 4154 16640 4160 16652
rect 3436 16612 4160 16640
rect 3436 16572 3464 16612
rect 4154 16600 4160 16612
rect 4212 16600 4218 16652
rect 5626 16640 5632 16652
rect 5539 16612 5632 16640
rect 5626 16600 5632 16612
rect 5684 16640 5690 16652
rect 7300 16640 7328 16736
rect 10042 16668 10048 16720
rect 10100 16708 10106 16720
rect 10100 16680 12664 16708
rect 10100 16668 10106 16680
rect 5684 16612 7328 16640
rect 5684 16600 5690 16612
rect 11514 16600 11520 16652
rect 11572 16640 11578 16652
rect 11793 16643 11851 16649
rect 11793 16640 11805 16643
rect 11572 16612 11805 16640
rect 11572 16600 11578 16612
rect 11793 16609 11805 16612
rect 11839 16609 11851 16643
rect 11793 16603 11851 16609
rect 12342 16600 12348 16652
rect 12400 16640 12406 16652
rect 12636 16649 12664 16680
rect 15010 16668 15016 16720
rect 15068 16708 15074 16720
rect 15764 16708 15792 16739
rect 15068 16680 15792 16708
rect 15068 16668 15074 16680
rect 12437 16643 12495 16649
rect 12437 16640 12449 16643
rect 12400 16612 12449 16640
rect 12400 16600 12406 16612
rect 12437 16609 12449 16612
rect 12483 16609 12495 16643
rect 12437 16603 12495 16609
rect 12621 16643 12679 16649
rect 12621 16609 12633 16643
rect 12667 16640 12679 16643
rect 12710 16640 12716 16652
rect 12667 16612 12716 16640
rect 12667 16609 12679 16612
rect 12621 16603 12679 16609
rect 12710 16600 12716 16612
rect 12768 16640 12774 16652
rect 13262 16640 13268 16652
rect 12768 16612 13268 16640
rect 12768 16600 12774 16612
rect 13262 16600 13268 16612
rect 13320 16600 13326 16652
rect 13446 16640 13452 16652
rect 13407 16612 13452 16640
rect 13446 16600 13452 16612
rect 13504 16600 13510 16652
rect 13725 16643 13783 16649
rect 13725 16609 13737 16643
rect 13771 16640 13783 16643
rect 13906 16640 13912 16652
rect 13771 16612 13912 16640
rect 13771 16609 13783 16612
rect 13725 16603 13783 16609
rect 13906 16600 13912 16612
rect 13964 16600 13970 16652
rect 14550 16600 14556 16652
rect 14608 16640 14614 16652
rect 14737 16643 14795 16649
rect 14737 16640 14749 16643
rect 14608 16612 14749 16640
rect 14608 16600 14614 16612
rect 14737 16609 14749 16612
rect 14783 16640 14795 16643
rect 14826 16640 14832 16652
rect 14783 16612 14832 16640
rect 14783 16609 14795 16612
rect 14737 16603 14795 16609
rect 14826 16600 14832 16612
rect 14884 16600 14890 16652
rect 14921 16643 14979 16649
rect 14921 16609 14933 16643
rect 14967 16609 14979 16643
rect 14921 16603 14979 16609
rect 15749 16643 15807 16649
rect 15749 16609 15761 16643
rect 15795 16640 15807 16643
rect 15856 16640 15884 16748
rect 17402 16736 17408 16748
rect 17460 16736 17466 16788
rect 20533 16779 20591 16785
rect 20533 16745 20545 16779
rect 20579 16776 20591 16779
rect 20990 16776 20996 16788
rect 20579 16748 20996 16776
rect 20579 16745 20591 16748
rect 20533 16739 20591 16745
rect 20990 16736 20996 16748
rect 21048 16736 21054 16788
rect 26510 16776 26516 16788
rect 25424 16748 26516 16776
rect 15948 16680 17264 16708
rect 15948 16649 15976 16680
rect 17236 16652 17264 16680
rect 17310 16668 17316 16720
rect 17368 16708 17374 16720
rect 18233 16711 18291 16717
rect 18233 16708 18245 16711
rect 17368 16680 18245 16708
rect 17368 16668 17374 16680
rect 18233 16677 18245 16680
rect 18279 16677 18291 16711
rect 21085 16711 21143 16717
rect 21085 16708 21097 16711
rect 18233 16671 18291 16677
rect 20548 16680 21097 16708
rect 15795 16612 15884 16640
rect 15933 16643 15991 16649
rect 15795 16609 15807 16612
rect 15749 16603 15807 16609
rect 15933 16609 15945 16643
rect 15979 16609 15991 16643
rect 16390 16640 16396 16652
rect 16351 16612 16396 16640
rect 15933 16603 15991 16609
rect 3160 16544 3464 16572
rect 6362 16532 6368 16584
rect 6420 16572 6426 16584
rect 6549 16575 6607 16581
rect 6549 16572 6561 16575
rect 6420 16544 6561 16572
rect 6420 16532 6426 16544
rect 6549 16541 6561 16544
rect 6595 16541 6607 16575
rect 6549 16535 6607 16541
rect 13538 16504 13544 16516
rect 13499 16476 13544 16504
rect 13538 16464 13544 16476
rect 13596 16464 13602 16516
rect 14936 16504 14964 16603
rect 16390 16600 16396 16612
rect 16448 16600 16454 16652
rect 16577 16643 16635 16649
rect 16577 16609 16589 16643
rect 16623 16609 16635 16643
rect 17218 16640 17224 16652
rect 17179 16612 17224 16640
rect 16577 16603 16635 16609
rect 16592 16572 16620 16603
rect 17218 16600 17224 16612
rect 17276 16600 17282 16652
rect 18598 16600 18604 16652
rect 18656 16640 18662 16652
rect 19061 16643 19119 16649
rect 19061 16640 19073 16643
rect 18656 16612 19073 16640
rect 18656 16600 18662 16612
rect 19061 16609 19073 16612
rect 19107 16640 19119 16643
rect 20257 16643 20315 16649
rect 19107 16612 19380 16640
rect 19107 16609 19119 16612
rect 19061 16603 19119 16609
rect 17310 16572 17316 16584
rect 16592 16544 17316 16572
rect 15470 16504 15476 16516
rect 14936 16476 15476 16504
rect 15470 16464 15476 16476
rect 15528 16504 15534 16516
rect 16592 16504 16620 16544
rect 17310 16532 17316 16544
rect 17368 16532 17374 16584
rect 15528 16476 16620 16504
rect 19352 16504 19380 16612
rect 20257 16609 20269 16643
rect 20303 16640 20315 16643
rect 20438 16640 20444 16652
rect 20303 16612 20444 16640
rect 20303 16609 20315 16612
rect 20257 16603 20315 16609
rect 20438 16600 20444 16612
rect 20496 16600 20502 16652
rect 20548 16581 20576 16680
rect 21085 16677 21097 16680
rect 21131 16677 21143 16711
rect 21085 16671 21143 16677
rect 20622 16600 20628 16652
rect 20680 16640 20686 16652
rect 20993 16643 21051 16649
rect 20993 16640 21005 16643
rect 20680 16612 21005 16640
rect 20680 16600 20686 16612
rect 20993 16609 21005 16612
rect 21039 16609 21051 16643
rect 20993 16603 21051 16609
rect 21177 16643 21235 16649
rect 21177 16609 21189 16643
rect 21223 16640 21235 16643
rect 22094 16640 22100 16652
rect 21223 16612 22100 16640
rect 21223 16609 21235 16612
rect 21177 16603 21235 16609
rect 22094 16600 22100 16612
rect 22152 16600 22158 16652
rect 23658 16640 23664 16652
rect 23400 16612 23664 16640
rect 20533 16575 20591 16581
rect 20533 16541 20545 16575
rect 20579 16541 20591 16575
rect 21082 16572 21088 16584
rect 20533 16535 20591 16541
rect 20640 16544 21088 16572
rect 20640 16504 20668 16544
rect 21082 16532 21088 16544
rect 21140 16572 21146 16584
rect 21910 16572 21916 16584
rect 21140 16544 21916 16572
rect 21140 16532 21146 16544
rect 21910 16532 21916 16544
rect 21968 16572 21974 16584
rect 23400 16572 23428 16612
rect 23658 16600 23664 16612
rect 23716 16600 23722 16652
rect 25222 16640 25228 16652
rect 25183 16612 25228 16640
rect 25222 16600 25228 16612
rect 25280 16600 25286 16652
rect 25424 16649 25452 16748
rect 26510 16736 26516 16748
rect 26568 16736 26574 16788
rect 32033 16779 32091 16785
rect 32033 16745 32045 16779
rect 32079 16776 32091 16779
rect 32122 16776 32128 16788
rect 32079 16748 32128 16776
rect 32079 16745 32091 16748
rect 32033 16739 32091 16745
rect 32122 16736 32128 16748
rect 32180 16736 32186 16788
rect 26973 16711 27031 16717
rect 25516 16680 26924 16708
rect 25409 16643 25467 16649
rect 25409 16609 25421 16643
rect 25455 16609 25467 16643
rect 25409 16603 25467 16609
rect 21968 16544 23428 16572
rect 25317 16575 25375 16581
rect 21968 16532 21974 16544
rect 25317 16541 25329 16575
rect 25363 16572 25375 16575
rect 25516 16572 25544 16680
rect 25682 16600 25688 16652
rect 25740 16640 25746 16652
rect 25961 16643 26019 16649
rect 25961 16640 25973 16643
rect 25740 16612 25973 16640
rect 25740 16600 25746 16612
rect 25961 16609 25973 16612
rect 26007 16609 26019 16643
rect 25961 16603 26019 16609
rect 26145 16643 26203 16649
rect 26145 16609 26157 16643
rect 26191 16609 26203 16643
rect 26145 16603 26203 16609
rect 25363 16544 25544 16572
rect 26160 16572 26188 16603
rect 26234 16600 26240 16652
rect 26292 16640 26298 16652
rect 26697 16643 26755 16649
rect 26697 16640 26709 16643
rect 26292 16612 26709 16640
rect 26292 16600 26298 16612
rect 26697 16609 26709 16612
rect 26743 16609 26755 16643
rect 26896 16640 26924 16680
rect 26973 16677 26985 16711
rect 27019 16708 27031 16711
rect 28534 16708 28540 16720
rect 27019 16680 28540 16708
rect 27019 16677 27031 16680
rect 26973 16671 27031 16677
rect 28534 16668 28540 16680
rect 28592 16668 28598 16720
rect 30834 16708 30840 16720
rect 30795 16680 30840 16708
rect 30834 16668 30840 16680
rect 30892 16668 30898 16720
rect 31938 16708 31944 16720
rect 31680 16680 31944 16708
rect 30558 16640 30564 16652
rect 26896 16612 27016 16640
rect 30519 16612 30564 16640
rect 26697 16603 26755 16609
rect 26418 16572 26424 16584
rect 26160 16544 26424 16572
rect 25363 16541 25375 16544
rect 25317 16535 25375 16541
rect 26418 16532 26424 16544
rect 26476 16532 26482 16584
rect 26988 16581 27016 16612
rect 30558 16600 30564 16612
rect 30616 16600 30622 16652
rect 30742 16600 30748 16652
rect 30800 16640 30806 16652
rect 31202 16640 31208 16652
rect 30800 16612 31208 16640
rect 30800 16600 30806 16612
rect 31202 16600 31208 16612
rect 31260 16600 31266 16652
rect 31386 16640 31392 16652
rect 31347 16612 31392 16640
rect 31386 16600 31392 16612
rect 31444 16600 31450 16652
rect 31570 16640 31576 16652
rect 31531 16612 31576 16640
rect 31570 16600 31576 16612
rect 31628 16600 31634 16652
rect 31680 16649 31708 16680
rect 31938 16668 31944 16680
rect 31996 16668 32002 16720
rect 32214 16668 32220 16720
rect 32272 16708 32278 16720
rect 32272 16680 32812 16708
rect 32272 16668 32278 16680
rect 31665 16643 31723 16649
rect 31665 16609 31677 16643
rect 31711 16609 31723 16643
rect 31665 16603 31723 16609
rect 31757 16643 31815 16649
rect 31757 16609 31769 16643
rect 31803 16640 31815 16643
rect 31846 16640 31852 16652
rect 31803 16612 31852 16640
rect 31803 16609 31815 16612
rect 31757 16603 31815 16609
rect 31846 16600 31852 16612
rect 31904 16640 31910 16652
rect 32784 16649 32812 16680
rect 32493 16643 32551 16649
rect 32493 16640 32505 16643
rect 31904 16612 32505 16640
rect 31904 16600 31910 16612
rect 32493 16609 32505 16612
rect 32539 16609 32551 16643
rect 32674 16643 32732 16649
rect 32674 16640 32686 16643
rect 32493 16603 32551 16609
rect 32600 16612 32686 16640
rect 26973 16575 27031 16581
rect 26973 16541 26985 16575
rect 27019 16541 27031 16575
rect 26973 16535 27031 16541
rect 32030 16532 32036 16584
rect 32088 16572 32094 16584
rect 32600 16572 32628 16612
rect 32674 16609 32686 16612
rect 32720 16609 32732 16643
rect 32674 16603 32732 16609
rect 32769 16643 32827 16649
rect 32769 16609 32781 16643
rect 32815 16609 32827 16643
rect 33413 16643 33471 16649
rect 33413 16640 33425 16643
rect 32769 16603 32827 16609
rect 32876 16612 33425 16640
rect 32876 16572 32904 16612
rect 33413 16609 33425 16612
rect 33459 16609 33471 16643
rect 33413 16603 33471 16609
rect 33502 16600 33508 16652
rect 33560 16640 33566 16652
rect 33560 16612 33605 16640
rect 33560 16600 33566 16612
rect 32088 16544 32904 16572
rect 32088 16532 32094 16544
rect 19352 16476 20668 16504
rect 15528 16464 15534 16476
rect 20806 16464 20812 16516
rect 20864 16504 20870 16516
rect 24762 16504 24768 16516
rect 20864 16476 24768 16504
rect 20864 16464 20870 16476
rect 24762 16464 24768 16476
rect 24820 16464 24826 16516
rect 26050 16464 26056 16516
rect 26108 16504 26114 16516
rect 26789 16507 26847 16513
rect 26789 16504 26801 16507
rect 26108 16476 26801 16504
rect 26108 16464 26114 16476
rect 26789 16473 26801 16476
rect 26835 16473 26847 16507
rect 26789 16467 26847 16473
rect 3050 16396 3056 16448
rect 3108 16436 3114 16448
rect 3329 16439 3387 16445
rect 3329 16436 3341 16439
rect 3108 16408 3341 16436
rect 3108 16396 3114 16408
rect 3329 16405 3341 16408
rect 3375 16405 3387 16439
rect 3329 16399 3387 16405
rect 15930 16396 15936 16448
rect 15988 16436 15994 16448
rect 16393 16439 16451 16445
rect 16393 16436 16405 16439
rect 15988 16408 16405 16436
rect 15988 16396 15994 16408
rect 16393 16405 16405 16408
rect 16439 16405 16451 16439
rect 16393 16399 16451 16405
rect 16942 16396 16948 16448
rect 17000 16436 17006 16448
rect 17129 16439 17187 16445
rect 17129 16436 17141 16439
rect 17000 16408 17141 16436
rect 17000 16396 17006 16408
rect 17129 16405 17141 16408
rect 17175 16405 17187 16439
rect 17129 16399 17187 16405
rect 19978 16396 19984 16448
rect 20036 16436 20042 16448
rect 20349 16439 20407 16445
rect 20349 16436 20361 16439
rect 20036 16408 20361 16436
rect 20036 16396 20042 16408
rect 20349 16405 20361 16408
rect 20395 16405 20407 16439
rect 20349 16399 20407 16405
rect 20438 16396 20444 16448
rect 20496 16436 20502 16448
rect 26145 16439 26203 16445
rect 26145 16436 26157 16439
rect 20496 16408 26157 16436
rect 20496 16396 20502 16408
rect 26145 16405 26157 16408
rect 26191 16436 26203 16439
rect 26510 16436 26516 16448
rect 26191 16408 26516 16436
rect 26191 16405 26203 16408
rect 26145 16399 26203 16405
rect 26510 16396 26516 16408
rect 26568 16396 26574 16448
rect 1104 16346 34316 16368
rect 1104 16294 6517 16346
rect 6569 16294 6581 16346
rect 6633 16294 6645 16346
rect 6697 16294 6709 16346
rect 6761 16294 17588 16346
rect 17640 16294 17652 16346
rect 17704 16294 17716 16346
rect 17768 16294 17780 16346
rect 17832 16294 28658 16346
rect 28710 16294 28722 16346
rect 28774 16294 28786 16346
rect 28838 16294 28850 16346
rect 28902 16294 34316 16346
rect 1104 16272 34316 16294
rect 4798 16232 4804 16244
rect 4759 16204 4804 16232
rect 4798 16192 4804 16204
rect 4856 16192 4862 16244
rect 14090 16232 14096 16244
rect 14051 16204 14096 16232
rect 14090 16192 14096 16204
rect 14148 16192 14154 16244
rect 14642 16192 14648 16244
rect 14700 16232 14706 16244
rect 15197 16235 15255 16241
rect 15197 16232 15209 16235
rect 14700 16204 15209 16232
rect 14700 16192 14706 16204
rect 15197 16201 15209 16204
rect 15243 16232 15255 16235
rect 16390 16232 16396 16244
rect 15243 16204 16396 16232
rect 15243 16201 15255 16204
rect 15197 16195 15255 16201
rect 16390 16192 16396 16204
rect 16448 16192 16454 16244
rect 18785 16235 18843 16241
rect 18785 16201 18797 16235
rect 18831 16232 18843 16235
rect 18966 16232 18972 16244
rect 18831 16204 18972 16232
rect 18831 16201 18843 16204
rect 18785 16195 18843 16201
rect 18966 16192 18972 16204
rect 19024 16192 19030 16244
rect 19518 16232 19524 16244
rect 19431 16204 19524 16232
rect 19518 16192 19524 16204
rect 19576 16232 19582 16244
rect 20622 16232 20628 16244
rect 19576 16204 20628 16232
rect 19576 16192 19582 16204
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 20898 16192 20904 16244
rect 20956 16232 20962 16244
rect 20956 16204 21220 16232
rect 20956 16192 20962 16204
rect 11149 16167 11207 16173
rect 11149 16133 11161 16167
rect 11195 16164 11207 16167
rect 11330 16164 11336 16176
rect 11195 16136 11336 16164
rect 11195 16133 11207 16136
rect 11149 16127 11207 16133
rect 11330 16124 11336 16136
rect 11388 16124 11394 16176
rect 12894 16164 12900 16176
rect 12820 16136 12900 16164
rect 3418 16096 3424 16108
rect 3379 16068 3424 16096
rect 3418 16056 3424 16068
rect 3476 16096 3482 16108
rect 9677 16099 9735 16105
rect 3476 16068 4476 16096
rect 3476 16056 3482 16068
rect 1394 16028 1400 16040
rect 1355 16000 1400 16028
rect 1394 15988 1400 16000
rect 1452 15988 1458 16040
rect 4154 16028 4160 16040
rect 4115 16000 4160 16028
rect 4154 15988 4160 16000
rect 4212 15988 4218 16040
rect 4448 16037 4476 16068
rect 9677 16065 9689 16099
rect 9723 16096 9735 16099
rect 10134 16096 10140 16108
rect 9723 16068 10140 16096
rect 9723 16065 9735 16068
rect 9677 16059 9735 16065
rect 10134 16056 10140 16068
rect 10192 16096 10198 16108
rect 10192 16068 11008 16096
rect 10192 16056 10198 16068
rect 4433 16031 4491 16037
rect 4433 15997 4445 16031
rect 4479 15997 4491 16031
rect 5166 16028 5172 16040
rect 5127 16000 5172 16028
rect 4433 15991 4491 15997
rect 5166 15988 5172 16000
rect 5224 15988 5230 16040
rect 6362 15988 6368 16040
rect 6420 16028 6426 16040
rect 6638 16028 6644 16040
rect 6420 16000 6644 16028
rect 6420 15988 6426 16000
rect 6638 15988 6644 16000
rect 6696 16028 6702 16040
rect 7285 16031 7343 16037
rect 7285 16028 7297 16031
rect 6696 16000 7297 16028
rect 6696 15988 6702 16000
rect 7285 15997 7297 16000
rect 7331 15997 7343 16031
rect 7285 15991 7343 15997
rect 9861 16031 9919 16037
rect 9861 15997 9873 16031
rect 9907 16028 9919 16031
rect 10870 16028 10876 16040
rect 9907 16000 10876 16028
rect 9907 15997 9919 16000
rect 9861 15991 9919 15997
rect 10870 15988 10876 16000
rect 10928 15988 10934 16040
rect 10980 16037 11008 16068
rect 10965 16031 11023 16037
rect 10965 15997 10977 16031
rect 11011 15997 11023 16031
rect 10965 15991 11023 15997
rect 12437 16031 12495 16037
rect 12437 15997 12449 16031
rect 12483 16028 12495 16031
rect 12820 16028 12848 16136
rect 12894 16124 12900 16136
rect 12952 16164 12958 16176
rect 16942 16164 16948 16176
rect 12952 16136 16948 16164
rect 12952 16124 12958 16136
rect 16942 16124 16948 16136
rect 17000 16124 17006 16176
rect 18877 16167 18935 16173
rect 18877 16133 18889 16167
rect 18923 16164 18935 16167
rect 19978 16164 19984 16176
rect 18923 16136 19984 16164
rect 18923 16133 18935 16136
rect 18877 16127 18935 16133
rect 19978 16124 19984 16136
rect 20036 16124 20042 16176
rect 13630 16096 13636 16108
rect 12912 16068 13636 16096
rect 12912 16037 12940 16068
rect 13630 16056 13636 16068
rect 13688 16056 13694 16108
rect 14826 16056 14832 16108
rect 14884 16096 14890 16108
rect 17126 16096 17132 16108
rect 14884 16068 17132 16096
rect 14884 16056 14890 16068
rect 12483 16000 12848 16028
rect 12897 16031 12955 16037
rect 12483 15997 12495 16000
rect 12437 15991 12495 15997
rect 12897 15997 12909 16031
rect 12943 15997 12955 16031
rect 12897 15991 12955 15997
rect 13354 15988 13360 16040
rect 13412 16028 13418 16040
rect 13909 16031 13967 16037
rect 13909 16028 13921 16031
rect 13412 16000 13921 16028
rect 13412 15988 13418 16000
rect 13909 15997 13921 16000
rect 13955 15997 13967 16031
rect 13909 15991 13967 15997
rect 14185 16031 14243 16037
rect 14185 15997 14197 16031
rect 14231 16028 14243 16031
rect 15930 16028 15936 16040
rect 14231 16000 15936 16028
rect 14231 15997 14243 16000
rect 14185 15991 14243 15997
rect 15930 15988 15936 16000
rect 15988 15988 15994 16040
rect 16040 16037 16068 16068
rect 17126 16056 17132 16068
rect 17184 16056 17190 16108
rect 18693 16099 18751 16105
rect 18693 16065 18705 16099
rect 18739 16096 18751 16099
rect 19794 16096 19800 16108
rect 18739 16068 19800 16096
rect 18739 16065 18751 16068
rect 18693 16059 18751 16065
rect 19794 16056 19800 16068
rect 19852 16056 19858 16108
rect 20990 16096 20996 16108
rect 20951 16068 20996 16096
rect 20990 16056 20996 16068
rect 21048 16056 21054 16108
rect 21192 16096 21220 16204
rect 22462 16192 22468 16244
rect 22520 16232 22526 16244
rect 22649 16235 22707 16241
rect 22649 16232 22661 16235
rect 22520 16204 22661 16232
rect 22520 16192 22526 16204
rect 22649 16201 22661 16204
rect 22695 16201 22707 16235
rect 26234 16232 26240 16244
rect 26195 16204 26240 16232
rect 22649 16195 22707 16201
rect 26234 16192 26240 16204
rect 26292 16192 26298 16244
rect 27893 16235 27951 16241
rect 27893 16201 27905 16235
rect 27939 16232 27951 16235
rect 28258 16232 28264 16244
rect 27939 16204 28264 16232
rect 27939 16201 27951 16204
rect 27893 16195 27951 16201
rect 26252 16164 26280 16192
rect 22572 16136 26280 16164
rect 21269 16099 21327 16105
rect 21269 16096 21281 16099
rect 21192 16068 21281 16096
rect 21269 16065 21281 16068
rect 21315 16096 21327 16099
rect 21726 16096 21732 16108
rect 21315 16068 21732 16096
rect 21315 16065 21327 16068
rect 21269 16059 21327 16065
rect 21726 16056 21732 16068
rect 21784 16056 21790 16108
rect 22572 16037 22600 16136
rect 22833 16099 22891 16105
rect 22833 16065 22845 16099
rect 22879 16096 22891 16099
rect 23385 16099 23443 16105
rect 23385 16096 23397 16099
rect 22879 16068 23397 16096
rect 22879 16065 22891 16068
rect 22833 16059 22891 16065
rect 23385 16065 23397 16068
rect 23431 16065 23443 16099
rect 23385 16059 23443 16065
rect 25222 16056 25228 16108
rect 25280 16096 25286 16108
rect 27908 16096 27936 16195
rect 28258 16192 28264 16204
rect 28316 16192 28322 16244
rect 29086 16192 29092 16244
rect 29144 16232 29150 16244
rect 30101 16235 30159 16241
rect 30101 16232 30113 16235
rect 29144 16204 30113 16232
rect 29144 16192 29150 16204
rect 30101 16201 30113 16204
rect 30147 16201 30159 16235
rect 30101 16195 30159 16201
rect 31018 16164 31024 16176
rect 25280 16068 27936 16096
rect 30484 16136 31024 16164
rect 25280 16056 25286 16068
rect 16025 16031 16083 16037
rect 16025 15997 16037 16031
rect 16071 15997 16083 16031
rect 16025 15991 16083 15997
rect 18969 16031 19027 16037
rect 18969 15997 18981 16031
rect 19015 16028 19027 16031
rect 22557 16031 22615 16037
rect 19015 16000 19748 16028
rect 19015 15997 19027 16000
rect 18969 15991 19027 15997
rect 1670 15960 1676 15972
rect 1631 15932 1676 15960
rect 1670 15920 1676 15932
rect 1728 15920 1734 15972
rect 2682 15920 2688 15972
rect 2740 15920 2746 15972
rect 7558 15960 7564 15972
rect 7519 15932 7564 15960
rect 7558 15920 7564 15932
rect 7616 15920 7622 15972
rect 8018 15920 8024 15972
rect 8076 15920 8082 15972
rect 8846 15920 8852 15972
rect 8904 15960 8910 15972
rect 11149 15963 11207 15969
rect 8904 15932 11100 15960
rect 8904 15920 8910 15932
rect 8202 15852 8208 15904
rect 8260 15892 8266 15904
rect 9033 15895 9091 15901
rect 9033 15892 9045 15895
rect 8260 15864 9045 15892
rect 8260 15852 8266 15864
rect 9033 15861 9045 15864
rect 9079 15861 9091 15895
rect 9033 15855 9091 15861
rect 10045 15895 10103 15901
rect 10045 15861 10057 15895
rect 10091 15892 10103 15895
rect 10870 15892 10876 15904
rect 10091 15864 10876 15892
rect 10091 15861 10103 15864
rect 10045 15855 10103 15861
rect 10870 15852 10876 15864
rect 10928 15852 10934 15904
rect 11072 15892 11100 15932
rect 11149 15929 11161 15963
rect 11195 15960 11207 15963
rect 15013 15963 15071 15969
rect 11195 15932 12434 15960
rect 11195 15929 11207 15932
rect 11149 15923 11207 15929
rect 12406 15904 12434 15932
rect 15013 15929 15025 15963
rect 15059 15929 15071 15963
rect 15013 15923 15071 15929
rect 15229 15963 15287 15969
rect 15229 15929 15241 15963
rect 15275 15960 15287 15963
rect 15746 15960 15752 15972
rect 15275 15932 15752 15960
rect 15275 15929 15287 15932
rect 15229 15923 15287 15929
rect 12253 15895 12311 15901
rect 12253 15892 12265 15895
rect 11072 15864 12265 15892
rect 12253 15861 12265 15864
rect 12299 15861 12311 15895
rect 12406 15864 12440 15904
rect 12253 15855 12311 15861
rect 12434 15852 12440 15864
rect 12492 15892 12498 15904
rect 12894 15892 12900 15904
rect 12492 15864 12900 15892
rect 12492 15852 12498 15864
rect 12894 15852 12900 15864
rect 12952 15852 12958 15904
rect 12989 15895 13047 15901
rect 12989 15861 13001 15895
rect 13035 15892 13047 15895
rect 13170 15892 13176 15904
rect 13035 15864 13176 15892
rect 13035 15861 13047 15864
rect 12989 15855 13047 15861
rect 13170 15852 13176 15864
rect 13228 15892 13234 15904
rect 13722 15892 13728 15904
rect 13228 15864 13728 15892
rect 13228 15852 13234 15864
rect 13722 15852 13728 15864
rect 13780 15852 13786 15904
rect 13906 15852 13912 15904
rect 13964 15892 13970 15904
rect 15028 15892 15056 15923
rect 15746 15920 15752 15932
rect 15804 15920 15810 15972
rect 17310 15920 17316 15972
rect 17368 15960 17374 15972
rect 19518 15960 19524 15972
rect 17368 15932 19524 15960
rect 17368 15920 17374 15932
rect 19518 15920 19524 15932
rect 19576 15920 19582 15972
rect 13964 15864 15056 15892
rect 15381 15895 15439 15901
rect 13964 15852 13970 15864
rect 15381 15861 15393 15895
rect 15427 15892 15439 15895
rect 15562 15892 15568 15904
rect 15427 15864 15568 15892
rect 15427 15861 15439 15864
rect 15381 15855 15439 15861
rect 15562 15852 15568 15864
rect 15620 15852 15626 15904
rect 15933 15895 15991 15901
rect 15933 15861 15945 15895
rect 15979 15892 15991 15895
rect 16206 15892 16212 15904
rect 15979 15864 16212 15892
rect 15979 15861 15991 15864
rect 15933 15855 15991 15861
rect 16206 15852 16212 15864
rect 16264 15852 16270 15904
rect 19720 15892 19748 16000
rect 22557 15997 22569 16031
rect 22603 15997 22615 16031
rect 22557 15991 22615 15997
rect 20530 15920 20536 15972
rect 20588 15920 20594 15972
rect 20714 15920 20720 15972
rect 20772 15960 20778 15972
rect 22572 15960 22600 15991
rect 23014 15988 23020 16040
rect 23072 16028 23078 16040
rect 23293 16031 23351 16037
rect 23293 16028 23305 16031
rect 23072 16000 23305 16028
rect 23072 15988 23078 16000
rect 23293 15997 23305 16000
rect 23339 15997 23351 16031
rect 23474 16028 23480 16040
rect 23435 16000 23480 16028
rect 23293 15991 23351 15997
rect 23474 15988 23480 16000
rect 23532 15988 23538 16040
rect 25501 16031 25559 16037
rect 25501 15997 25513 16031
rect 25547 16028 25559 16031
rect 25590 16028 25596 16040
rect 25547 16000 25596 16028
rect 25547 15997 25559 16000
rect 25501 15991 25559 15997
rect 25590 15988 25596 16000
rect 25648 15988 25654 16040
rect 25700 16037 25728 16068
rect 25685 16031 25743 16037
rect 25685 15997 25697 16031
rect 25731 15997 25743 16031
rect 25685 15991 25743 15997
rect 26145 16031 26203 16037
rect 26145 15997 26157 16031
rect 26191 15997 26203 16031
rect 26326 16028 26332 16040
rect 26287 16000 26332 16028
rect 26145 15991 26203 15997
rect 20772 15932 22600 15960
rect 20772 15920 20778 15932
rect 22738 15920 22744 15972
rect 22796 15960 22802 15972
rect 25314 15960 25320 15972
rect 22796 15932 25320 15960
rect 22796 15920 22802 15932
rect 25314 15920 25320 15932
rect 25372 15920 25378 15972
rect 25608 15960 25636 15988
rect 26160 15960 26188 15991
rect 26326 15988 26332 16000
rect 26384 15988 26390 16040
rect 28534 15988 28540 16040
rect 28592 16028 28598 16040
rect 29006 16031 29064 16037
rect 29006 16028 29018 16031
rect 28592 16000 29018 16028
rect 28592 15988 28598 16000
rect 29006 15997 29018 16000
rect 29052 15997 29064 16031
rect 29006 15991 29064 15997
rect 29178 15988 29184 16040
rect 29236 16028 29242 16040
rect 30484 16037 30512 16136
rect 31018 16124 31024 16136
rect 31076 16124 31082 16176
rect 31570 16096 31576 16108
rect 30668 16068 31576 16096
rect 30668 16040 30696 16068
rect 31570 16056 31576 16068
rect 31628 16056 31634 16108
rect 29273 16031 29331 16037
rect 29273 16028 29285 16031
rect 29236 16000 29285 16028
rect 29236 15988 29242 16000
rect 29273 15997 29285 16000
rect 29319 15997 29331 16031
rect 29273 15991 29331 15997
rect 30377 16031 30435 16037
rect 30377 15997 30389 16031
rect 30423 15997 30435 16031
rect 30377 15991 30435 15997
rect 30466 16031 30524 16037
rect 30466 15997 30478 16031
rect 30512 15997 30524 16031
rect 30466 15991 30524 15997
rect 30561 16031 30619 16037
rect 30561 15997 30573 16031
rect 30607 16028 30619 16031
rect 30650 16028 30656 16040
rect 30607 16000 30656 16028
rect 30607 15997 30619 16000
rect 30561 15991 30619 15997
rect 25608 15932 26188 15960
rect 30392 15960 30420 15991
rect 30650 15988 30656 16000
rect 30708 15988 30714 16040
rect 30745 16031 30803 16037
rect 30745 15997 30757 16031
rect 30791 16028 30803 16031
rect 31386 16028 31392 16040
rect 30791 16000 31392 16028
rect 30791 15997 30803 16000
rect 30745 15991 30803 15997
rect 31386 15988 31392 16000
rect 31444 15988 31450 16040
rect 31757 16031 31815 16037
rect 31757 15997 31769 16031
rect 31803 16028 31815 16031
rect 31846 16028 31852 16040
rect 31803 16000 31852 16028
rect 31803 15997 31815 16000
rect 31757 15991 31815 15997
rect 31846 15988 31852 16000
rect 31904 15988 31910 16040
rect 33594 16028 33600 16040
rect 33555 16000 33600 16028
rect 33594 15988 33600 16000
rect 33652 15988 33658 16040
rect 30834 15960 30840 15972
rect 30392 15932 30840 15960
rect 30834 15920 30840 15932
rect 30892 15920 30898 15972
rect 31202 15920 31208 15972
rect 31260 15960 31266 15972
rect 31941 15963 31999 15969
rect 31941 15960 31953 15963
rect 31260 15932 31953 15960
rect 31260 15920 31266 15932
rect 31941 15929 31953 15932
rect 31987 15960 31999 15963
rect 33505 15963 33563 15969
rect 33505 15960 33517 15963
rect 31987 15932 33517 15960
rect 31987 15929 31999 15932
rect 31941 15923 31999 15929
rect 33505 15929 33517 15932
rect 33551 15929 33563 15963
rect 33505 15923 33563 15929
rect 20806 15892 20812 15904
rect 19720 15864 20812 15892
rect 20806 15852 20812 15864
rect 20864 15852 20870 15904
rect 22002 15852 22008 15904
rect 22060 15892 22066 15904
rect 22833 15895 22891 15901
rect 22833 15892 22845 15895
rect 22060 15864 22845 15892
rect 22060 15852 22066 15864
rect 22833 15861 22845 15864
rect 22879 15861 22891 15895
rect 32122 15892 32128 15904
rect 32083 15864 32128 15892
rect 22833 15855 22891 15861
rect 32122 15852 32128 15864
rect 32180 15852 32186 15904
rect 1104 15802 34316 15824
rect 1104 15750 12052 15802
rect 12104 15750 12116 15802
rect 12168 15750 12180 15802
rect 12232 15750 12244 15802
rect 12296 15750 23123 15802
rect 23175 15750 23187 15802
rect 23239 15750 23251 15802
rect 23303 15750 23315 15802
rect 23367 15750 34316 15802
rect 1104 15728 34316 15750
rect 1670 15648 1676 15700
rect 1728 15688 1734 15700
rect 2869 15691 2927 15697
rect 2869 15688 2881 15691
rect 1728 15660 2881 15688
rect 1728 15648 1734 15660
rect 2869 15657 2881 15660
rect 2915 15657 2927 15691
rect 7006 15688 7012 15700
rect 2869 15651 2927 15657
rect 5184 15660 7012 15688
rect 2682 15580 2688 15632
rect 2740 15620 2746 15632
rect 5184 15620 5212 15660
rect 7006 15648 7012 15660
rect 7064 15688 7070 15700
rect 8018 15688 8024 15700
rect 7064 15660 8024 15688
rect 7064 15648 7070 15660
rect 8018 15648 8024 15660
rect 8076 15688 8082 15700
rect 9766 15688 9772 15700
rect 8076 15660 9772 15688
rect 8076 15648 8082 15660
rect 9766 15648 9772 15660
rect 9824 15688 9830 15700
rect 9824 15660 10456 15688
rect 9824 15648 9830 15660
rect 2740 15606 5212 15620
rect 2740 15592 5198 15606
rect 2740 15580 2746 15592
rect 7282 15580 7288 15632
rect 7340 15620 7346 15632
rect 7466 15620 7472 15632
rect 7340 15592 7472 15620
rect 7340 15580 7346 15592
rect 7466 15580 7472 15592
rect 7524 15620 7530 15632
rect 8481 15623 8539 15629
rect 8481 15620 8493 15623
rect 7524 15592 8493 15620
rect 7524 15580 7530 15592
rect 8481 15589 8493 15592
rect 8527 15589 8539 15623
rect 9674 15620 9680 15632
rect 9635 15592 9680 15620
rect 8481 15583 8539 15589
rect 9674 15580 9680 15592
rect 9732 15580 9738 15632
rect 10428 15629 10456 15660
rect 15378 15648 15384 15700
rect 15436 15688 15442 15700
rect 16393 15691 16451 15697
rect 16393 15688 16405 15691
rect 15436 15660 16405 15688
rect 15436 15648 15442 15660
rect 16393 15657 16405 15660
rect 16439 15688 16451 15691
rect 16439 15660 17448 15688
rect 16439 15657 16451 15660
rect 16393 15651 16451 15657
rect 10413 15623 10471 15629
rect 10413 15589 10425 15623
rect 10459 15620 10471 15623
rect 10962 15620 10968 15632
rect 10459 15592 10968 15620
rect 10459 15589 10471 15592
rect 10413 15583 10471 15589
rect 10962 15580 10968 15592
rect 11020 15580 11026 15632
rect 13078 15620 13084 15632
rect 12636 15592 13084 15620
rect 3050 15552 3056 15564
rect 3011 15524 3056 15552
rect 3050 15512 3056 15524
rect 3108 15512 3114 15564
rect 3329 15555 3387 15561
rect 3329 15521 3341 15555
rect 3375 15552 3387 15555
rect 3418 15552 3424 15564
rect 3375 15524 3424 15552
rect 3375 15521 3387 15524
rect 3329 15515 3387 15521
rect 3418 15512 3424 15524
rect 3476 15512 3482 15564
rect 7653 15555 7711 15561
rect 7653 15521 7665 15555
rect 7699 15552 7711 15555
rect 8202 15552 8208 15564
rect 7699 15524 8208 15552
rect 7699 15521 7711 15524
rect 7653 15515 7711 15521
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 10870 15512 10876 15564
rect 10928 15552 10934 15564
rect 11057 15555 11115 15561
rect 11057 15552 11069 15555
rect 10928 15524 11069 15552
rect 10928 15512 10934 15524
rect 11057 15521 11069 15524
rect 11103 15521 11115 15555
rect 11057 15515 11115 15521
rect 11149 15555 11207 15561
rect 11149 15521 11161 15555
rect 11195 15521 11207 15555
rect 11149 15515 11207 15521
rect 2958 15444 2964 15496
rect 3016 15484 3022 15496
rect 3237 15487 3295 15493
rect 3237 15484 3249 15487
rect 3016 15456 3249 15484
rect 3016 15444 3022 15456
rect 3237 15453 3249 15456
rect 3283 15484 3295 15487
rect 4062 15484 4068 15496
rect 3283 15456 4068 15484
rect 3283 15453 3295 15456
rect 3237 15447 3295 15453
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 6362 15484 6368 15496
rect 6323 15456 6368 15484
rect 6362 15444 6368 15456
rect 6420 15444 6426 15496
rect 6638 15484 6644 15496
rect 6551 15456 6644 15484
rect 6638 15444 6644 15456
rect 6696 15444 6702 15496
rect 7834 15484 7840 15496
rect 7795 15456 7840 15484
rect 7834 15444 7840 15456
rect 7892 15444 7898 15496
rect 4522 15308 4528 15360
rect 4580 15348 4586 15360
rect 4893 15351 4951 15357
rect 4893 15348 4905 15351
rect 4580 15320 4905 15348
rect 4580 15308 4586 15320
rect 4893 15317 4905 15320
rect 4939 15348 4951 15351
rect 5166 15348 5172 15360
rect 4939 15320 5172 15348
rect 4939 15317 4951 15320
rect 4893 15311 4951 15317
rect 5166 15308 5172 15320
rect 5224 15308 5230 15360
rect 5994 15308 6000 15360
rect 6052 15348 6058 15360
rect 6656 15348 6684 15444
rect 8294 15416 8300 15428
rect 8255 15388 8300 15416
rect 8294 15376 8300 15388
rect 8352 15376 8358 15428
rect 11164 15416 11192 15515
rect 11238 15512 11244 15564
rect 11296 15552 11302 15564
rect 11425 15555 11483 15561
rect 11425 15552 11437 15555
rect 11296 15524 11437 15552
rect 11296 15512 11302 15524
rect 11425 15521 11437 15524
rect 11471 15521 11483 15555
rect 11425 15515 11483 15521
rect 11330 15484 11336 15496
rect 11291 15456 11336 15484
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 12636 15493 12664 15592
rect 13078 15580 13084 15592
rect 13136 15580 13142 15632
rect 17310 15620 17316 15632
rect 17271 15592 17316 15620
rect 17310 15580 17316 15592
rect 17368 15580 17374 15632
rect 12805 15555 12863 15561
rect 12805 15521 12817 15555
rect 12851 15552 12863 15555
rect 12894 15552 12900 15564
rect 12851 15524 12900 15552
rect 12851 15521 12863 15524
rect 12805 15515 12863 15521
rect 12894 15512 12900 15524
rect 12952 15512 12958 15564
rect 13354 15512 13360 15564
rect 13412 15552 13418 15564
rect 13633 15555 13691 15561
rect 13633 15552 13645 15555
rect 13412 15524 13645 15552
rect 13412 15512 13418 15524
rect 13633 15521 13645 15524
rect 13679 15521 13691 15555
rect 13633 15515 13691 15521
rect 13722 15512 13728 15564
rect 13780 15552 13786 15564
rect 15381 15555 15439 15561
rect 15381 15552 15393 15555
rect 13780 15524 15393 15552
rect 13780 15512 13786 15524
rect 15381 15521 15393 15524
rect 15427 15521 15439 15555
rect 15562 15552 15568 15564
rect 15523 15524 15568 15552
rect 15381 15515 15439 15521
rect 15562 15512 15568 15524
rect 15620 15552 15626 15564
rect 16209 15555 16267 15561
rect 16209 15552 16221 15555
rect 15620 15524 16221 15552
rect 15620 15512 15626 15524
rect 16209 15521 16221 15524
rect 16255 15521 16267 15555
rect 16209 15515 16267 15521
rect 16574 15512 16580 15564
rect 16632 15552 16638 15564
rect 17083 15555 17141 15561
rect 17083 15552 17095 15555
rect 16632 15524 17095 15552
rect 16632 15512 16638 15524
rect 17083 15521 17095 15524
rect 17129 15521 17141 15555
rect 17218 15552 17224 15564
rect 17179 15524 17224 15552
rect 17083 15515 17141 15521
rect 17218 15512 17224 15524
rect 17276 15512 17282 15564
rect 17420 15561 17448 15660
rect 20530 15648 20536 15700
rect 20588 15688 20594 15700
rect 20714 15688 20720 15700
rect 20588 15660 20720 15688
rect 20588 15648 20594 15660
rect 20714 15648 20720 15660
rect 20772 15688 20778 15700
rect 21910 15688 21916 15700
rect 20772 15660 21916 15688
rect 20772 15648 20778 15660
rect 21910 15648 21916 15660
rect 21968 15688 21974 15700
rect 23474 15688 23480 15700
rect 21968 15660 22508 15688
rect 23435 15660 23480 15688
rect 21968 15648 21974 15660
rect 22002 15620 22008 15632
rect 21963 15592 22008 15620
rect 22002 15580 22008 15592
rect 22060 15580 22066 15632
rect 22480 15606 22508 15660
rect 23474 15648 23480 15660
rect 23532 15648 23538 15700
rect 30834 15648 30840 15700
rect 30892 15688 30898 15700
rect 32030 15688 32036 15700
rect 30892 15660 31432 15688
rect 30892 15648 30898 15660
rect 17405 15555 17463 15561
rect 17405 15521 17417 15555
rect 17451 15552 17463 15555
rect 17862 15552 17868 15564
rect 17451 15524 17868 15552
rect 17451 15521 17463 15524
rect 17405 15515 17463 15521
rect 17862 15512 17868 15524
rect 17920 15512 17926 15564
rect 21726 15552 21732 15564
rect 21687 15524 21732 15552
rect 21726 15512 21732 15524
rect 21784 15512 21790 15564
rect 23492 15552 23520 15648
rect 25866 15620 25872 15632
rect 25516 15592 25872 15620
rect 25516 15561 25544 15592
rect 25866 15580 25872 15592
rect 25924 15620 25930 15632
rect 26050 15620 26056 15632
rect 25924 15592 26056 15620
rect 25924 15580 25930 15592
rect 26050 15580 26056 15592
rect 26108 15580 26114 15632
rect 27982 15620 27988 15632
rect 26160 15592 27988 15620
rect 23937 15555 23995 15561
rect 23937 15552 23949 15555
rect 23492 15524 23949 15552
rect 23937 15521 23949 15524
rect 23983 15521 23995 15555
rect 23937 15515 23995 15521
rect 25501 15555 25559 15561
rect 25501 15521 25513 15555
rect 25547 15521 25559 15555
rect 25501 15515 25559 15521
rect 25682 15512 25688 15564
rect 25740 15552 25746 15564
rect 26160 15561 26188 15592
rect 27982 15580 27988 15592
rect 28040 15580 28046 15632
rect 31404 15629 31432 15660
rect 31772 15660 32036 15688
rect 31205 15623 31263 15629
rect 31205 15589 31217 15623
rect 31251 15589 31263 15623
rect 31205 15583 31263 15589
rect 31389 15623 31447 15629
rect 31389 15589 31401 15623
rect 31435 15589 31447 15623
rect 31389 15583 31447 15589
rect 25961 15555 26019 15561
rect 25961 15552 25973 15555
rect 25740 15524 25973 15552
rect 25740 15512 25746 15524
rect 25961 15521 25973 15524
rect 26007 15521 26019 15555
rect 25961 15515 26019 15521
rect 26145 15555 26203 15561
rect 26145 15521 26157 15555
rect 26191 15521 26203 15555
rect 26145 15515 26203 15521
rect 26602 15512 26608 15564
rect 26660 15552 26666 15564
rect 26789 15555 26847 15561
rect 26789 15552 26801 15555
rect 26660 15524 26801 15552
rect 26660 15512 26666 15524
rect 26789 15521 26801 15524
rect 26835 15521 26847 15555
rect 26789 15515 26847 15521
rect 26973 15555 27031 15561
rect 26973 15521 26985 15555
rect 27019 15521 27031 15555
rect 26973 15515 27031 15521
rect 12529 15487 12587 15493
rect 12529 15453 12541 15487
rect 12575 15453 12587 15487
rect 12529 15447 12587 15453
rect 12621 15487 12679 15493
rect 12621 15453 12633 15487
rect 12667 15453 12679 15487
rect 12621 15447 12679 15453
rect 12713 15487 12771 15493
rect 12713 15453 12725 15487
rect 12759 15484 12771 15487
rect 13446 15484 13452 15496
rect 12759 15456 13452 15484
rect 12759 15453 12771 15456
rect 12713 15447 12771 15453
rect 12345 15419 12403 15425
rect 12345 15416 12357 15419
rect 11164 15388 12357 15416
rect 12345 15385 12357 15388
rect 12391 15385 12403 15419
rect 12544 15416 12572 15447
rect 13446 15444 13452 15456
rect 13504 15444 13510 15496
rect 15289 15487 15347 15493
rect 15289 15453 15301 15487
rect 15335 15484 15347 15487
rect 16666 15484 16672 15496
rect 15335 15456 16672 15484
rect 15335 15453 15347 15456
rect 15289 15447 15347 15453
rect 16666 15444 16672 15456
rect 16724 15444 16730 15496
rect 16945 15487 17003 15493
rect 16945 15453 16957 15487
rect 16991 15484 17003 15487
rect 19058 15484 19064 15496
rect 16991 15456 19064 15484
rect 16991 15453 17003 15456
rect 16945 15447 17003 15453
rect 19058 15444 19064 15456
rect 19116 15444 19122 15496
rect 25222 15484 25228 15496
rect 25183 15456 25228 15484
rect 25222 15444 25228 15456
rect 25280 15444 25286 15496
rect 26326 15444 26332 15496
rect 26384 15484 26390 15496
rect 26988 15484 27016 15515
rect 27706 15512 27712 15564
rect 27764 15552 27770 15564
rect 27873 15555 27931 15561
rect 27873 15552 27885 15555
rect 27764 15524 27885 15552
rect 27764 15512 27770 15524
rect 27873 15521 27885 15524
rect 27919 15521 27931 15555
rect 31220 15552 31248 15583
rect 31772 15552 31800 15660
rect 32030 15648 32036 15660
rect 32088 15648 32094 15700
rect 33594 15688 33600 15700
rect 33555 15660 33600 15688
rect 33594 15648 33600 15660
rect 33652 15648 33658 15700
rect 31846 15580 31852 15632
rect 31904 15620 31910 15632
rect 32125 15623 32183 15629
rect 32125 15620 32137 15623
rect 31904 15592 32137 15620
rect 31904 15580 31910 15592
rect 32125 15589 32137 15592
rect 32171 15589 32183 15623
rect 32125 15583 32183 15589
rect 32582 15580 32588 15632
rect 32640 15580 32646 15632
rect 31220 15524 31800 15552
rect 27873 15515 27931 15521
rect 27614 15484 27620 15496
rect 26384 15456 27016 15484
rect 27575 15456 27620 15484
rect 26384 15444 26390 15456
rect 12802 15416 12808 15428
rect 12544 15388 12808 15416
rect 12345 15379 12403 15385
rect 12802 15376 12808 15388
rect 12860 15376 12866 15428
rect 7466 15348 7472 15360
rect 6052 15320 6684 15348
rect 7427 15320 7472 15348
rect 6052 15308 6058 15320
rect 7466 15308 7472 15320
rect 7524 15308 7530 15360
rect 10502 15308 10508 15360
rect 10560 15348 10566 15360
rect 10873 15351 10931 15357
rect 10873 15348 10885 15351
rect 10560 15320 10885 15348
rect 10560 15308 10566 15320
rect 10873 15317 10885 15320
rect 10919 15317 10931 15351
rect 10873 15311 10931 15317
rect 11790 15308 11796 15360
rect 11848 15348 11854 15360
rect 12710 15348 12716 15360
rect 11848 15320 12716 15348
rect 11848 15308 11854 15320
rect 12710 15308 12716 15320
rect 12768 15348 12774 15360
rect 13449 15351 13507 15357
rect 13449 15348 13461 15351
rect 12768 15320 13461 15348
rect 12768 15308 12774 15320
rect 13449 15317 13461 15320
rect 13495 15317 13507 15351
rect 15746 15348 15752 15360
rect 15707 15320 15752 15348
rect 13449 15311 13507 15317
rect 15746 15308 15752 15320
rect 15804 15308 15810 15360
rect 17402 15308 17408 15360
rect 17460 15348 17466 15360
rect 17589 15351 17647 15357
rect 17589 15348 17601 15351
rect 17460 15320 17601 15348
rect 17460 15308 17466 15320
rect 17589 15317 17601 15320
rect 17635 15317 17647 15351
rect 17589 15311 17647 15317
rect 23934 15308 23940 15360
rect 23992 15348 23998 15360
rect 24029 15351 24087 15357
rect 24029 15348 24041 15351
rect 23992 15320 24041 15348
rect 23992 15308 23998 15320
rect 24029 15317 24041 15320
rect 24075 15317 24087 15351
rect 25314 15348 25320 15360
rect 25275 15320 25320 15348
rect 24029 15311 24087 15317
rect 25314 15308 25320 15320
rect 25372 15308 25378 15360
rect 25409 15351 25467 15357
rect 25409 15317 25421 15351
rect 25455 15348 25467 15351
rect 26050 15348 26056 15360
rect 25455 15320 26056 15348
rect 25455 15317 25467 15320
rect 25409 15311 25467 15317
rect 26050 15308 26056 15320
rect 26108 15308 26114 15360
rect 26786 15308 26792 15360
rect 26844 15348 26850 15360
rect 26881 15351 26939 15357
rect 26881 15348 26893 15351
rect 26844 15320 26893 15348
rect 26844 15308 26850 15320
rect 26881 15317 26893 15320
rect 26927 15317 26939 15351
rect 26988 15348 27016 15456
rect 27614 15444 27620 15456
rect 27672 15444 27678 15496
rect 31754 15444 31760 15496
rect 31812 15484 31818 15496
rect 31849 15487 31907 15493
rect 31849 15484 31861 15487
rect 31812 15456 31861 15484
rect 31812 15444 31818 15456
rect 31849 15453 31861 15456
rect 31895 15453 31907 15487
rect 31849 15447 31907 15453
rect 28997 15351 29055 15357
rect 28997 15348 29009 15351
rect 26988 15320 29009 15348
rect 26881 15311 26939 15317
rect 28997 15317 29009 15320
rect 29043 15317 29055 15351
rect 31018 15348 31024 15360
rect 30979 15320 31024 15348
rect 28997 15311 29055 15317
rect 31018 15308 31024 15320
rect 31076 15308 31082 15360
rect 31202 15348 31208 15360
rect 31163 15320 31208 15348
rect 31202 15308 31208 15320
rect 31260 15308 31266 15360
rect 1104 15258 34316 15280
rect 1104 15206 6517 15258
rect 6569 15206 6581 15258
rect 6633 15206 6645 15258
rect 6697 15206 6709 15258
rect 6761 15206 17588 15258
rect 17640 15206 17652 15258
rect 17704 15206 17716 15258
rect 17768 15206 17780 15258
rect 17832 15206 28658 15258
rect 28710 15206 28722 15258
rect 28774 15206 28786 15258
rect 28838 15206 28850 15258
rect 28902 15206 34316 15258
rect 1104 15184 34316 15206
rect 10042 15104 10048 15156
rect 10100 15144 10106 15156
rect 12161 15147 12219 15153
rect 12161 15144 12173 15147
rect 10100 15116 12173 15144
rect 10100 15104 10106 15116
rect 12161 15113 12173 15116
rect 12207 15113 12219 15147
rect 13173 15147 13231 15153
rect 13173 15144 13185 15147
rect 12161 15107 12219 15113
rect 12406 15116 13185 15144
rect 3418 15036 3424 15088
rect 3476 15076 3482 15088
rect 3476 15048 4752 15076
rect 3476 15036 3482 15048
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 3973 15011 4031 15017
rect 3973 15008 3985 15011
rect 1719 14980 3985 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 3973 14977 3985 14980
rect 4019 14977 4031 15011
rect 3973 14971 4031 14977
rect 4062 14968 4068 15020
rect 4120 15008 4126 15020
rect 4724 15017 4752 15048
rect 11054 15036 11060 15088
rect 11112 15076 11118 15088
rect 12406 15076 12434 15116
rect 13173 15113 13185 15116
rect 13219 15113 13231 15147
rect 13173 15107 13231 15113
rect 17402 15104 17408 15156
rect 17460 15104 17466 15156
rect 17954 15104 17960 15156
rect 18012 15144 18018 15156
rect 21818 15144 21824 15156
rect 18012 15116 21824 15144
rect 18012 15104 18018 15116
rect 21818 15104 21824 15116
rect 21876 15104 21882 15156
rect 24946 15144 24952 15156
rect 24228 15116 24952 15144
rect 11112 15048 12434 15076
rect 11112 15036 11118 15048
rect 4709 15011 4767 15017
rect 4120 14980 4165 15008
rect 4120 14968 4126 14980
rect 4709 14977 4721 15011
rect 4755 15008 4767 15011
rect 5074 15008 5080 15020
rect 4755 14980 5080 15008
rect 4755 14977 4767 14980
rect 4709 14971 4767 14977
rect 5074 14968 5080 14980
rect 5132 15008 5138 15020
rect 5445 15011 5503 15017
rect 5445 15008 5457 15011
rect 5132 14980 5457 15008
rect 5132 14968 5138 14980
rect 5445 14977 5457 14980
rect 5491 14977 5503 15011
rect 10502 15008 10508 15020
rect 10463 14980 10508 15008
rect 5445 14971 5503 14977
rect 10502 14968 10508 14980
rect 10560 14968 10566 15020
rect 10778 15008 10784 15020
rect 10739 14980 10784 15008
rect 10778 14968 10784 14980
rect 10836 14968 10842 15020
rect 13630 14968 13636 15020
rect 13688 15008 13694 15020
rect 14553 15011 14611 15017
rect 14553 15008 14565 15011
rect 13688 14980 14565 15008
rect 13688 14968 13694 14980
rect 14553 14977 14565 14980
rect 14599 14977 14611 15011
rect 16390 15008 16396 15020
rect 14553 14971 14611 14977
rect 15488 14980 16396 15008
rect 15488 14952 15516 14980
rect 16390 14968 16396 14980
rect 16448 14968 16454 15020
rect 17420 15008 17448 15104
rect 20717 15079 20775 15085
rect 20717 15045 20729 15079
rect 20763 15076 20775 15079
rect 22462 15076 22468 15088
rect 20763 15048 22468 15076
rect 20763 15045 20775 15048
rect 20717 15039 20775 15045
rect 22462 15036 22468 15048
rect 22520 15036 22526 15088
rect 17589 15011 17647 15017
rect 17589 15008 17601 15011
rect 17420 14980 17601 15008
rect 17589 14977 17601 14980
rect 17635 14977 17647 15011
rect 17589 14971 17647 14977
rect 20901 15011 20959 15017
rect 20901 14977 20913 15011
rect 20947 15008 20959 15011
rect 22278 15008 22284 15020
rect 20947 14980 22284 15008
rect 20947 14977 20959 14980
rect 20901 14971 20959 14977
rect 22278 14968 22284 14980
rect 22336 14968 22342 15020
rect 24228 15017 24256 15116
rect 24946 15104 24952 15116
rect 25004 15104 25010 15156
rect 25593 15147 25651 15153
rect 25593 15113 25605 15147
rect 25639 15144 25651 15147
rect 25774 15144 25780 15156
rect 25639 15116 25780 15144
rect 25639 15113 25651 15116
rect 25593 15107 25651 15113
rect 25774 15104 25780 15116
rect 25832 15104 25838 15156
rect 25866 15104 25872 15156
rect 25924 15144 25930 15156
rect 26605 15147 26663 15153
rect 26605 15144 26617 15147
rect 25924 15116 26617 15144
rect 25924 15104 25930 15116
rect 26605 15113 26617 15116
rect 26651 15113 26663 15147
rect 26605 15107 26663 15113
rect 26697 15147 26755 15153
rect 26697 15113 26709 15147
rect 26743 15144 26755 15147
rect 27706 15144 27712 15156
rect 26743 15116 27712 15144
rect 26743 15113 26755 15116
rect 26697 15107 26755 15113
rect 27706 15104 27712 15116
rect 27764 15104 27770 15156
rect 30742 15144 30748 15156
rect 30703 15116 30748 15144
rect 30742 15104 30748 15116
rect 30800 15104 30806 15156
rect 31846 15144 31852 15156
rect 31807 15116 31852 15144
rect 31846 15104 31852 15116
rect 31904 15104 31910 15156
rect 24213 15011 24271 15017
rect 24213 14977 24225 15011
rect 24259 14977 24271 15011
rect 26786 15008 26792 15020
rect 26747 14980 26792 15008
rect 24213 14971 24271 14977
rect 26786 14968 26792 14980
rect 26844 14968 26850 15020
rect 27614 14968 27620 15020
rect 27672 15008 27678 15020
rect 28994 15008 29000 15020
rect 27672 14980 29000 15008
rect 27672 14968 27678 14980
rect 28994 14968 29000 14980
rect 29052 15008 29058 15020
rect 31662 15008 31668 15020
rect 29052 14980 31668 15008
rect 29052 14968 29058 14980
rect 31662 14968 31668 14980
rect 31720 14968 31726 15020
rect 1394 14940 1400 14952
rect 1355 14912 1400 14940
rect 1394 14900 1400 14912
rect 1452 14900 1458 14952
rect 3326 14900 3332 14952
rect 3384 14940 3390 14952
rect 3881 14943 3939 14949
rect 3881 14940 3893 14943
rect 3384 14912 3893 14940
rect 3384 14900 3390 14912
rect 3881 14909 3893 14912
rect 3927 14909 3939 14943
rect 3881 14903 3939 14909
rect 4246 14900 4252 14952
rect 4304 14940 4310 14952
rect 4341 14943 4399 14949
rect 4341 14940 4353 14943
rect 4304 14912 4353 14940
rect 4304 14900 4310 14912
rect 4341 14909 4353 14912
rect 4387 14940 4399 14943
rect 5166 14940 5172 14952
rect 4387 14912 5172 14940
rect 4387 14909 4399 14912
rect 4341 14903 4399 14909
rect 5166 14900 5172 14912
rect 5224 14900 5230 14952
rect 5537 14943 5595 14949
rect 5537 14909 5549 14943
rect 5583 14909 5595 14943
rect 7834 14940 7840 14952
rect 7795 14912 7840 14940
rect 5537 14903 5595 14909
rect 2682 14832 2688 14884
rect 2740 14832 2746 14884
rect 3421 14875 3479 14881
rect 3421 14841 3433 14875
rect 3467 14872 3479 14875
rect 4154 14872 4160 14884
rect 3467 14844 4160 14872
rect 3467 14841 3479 14844
rect 3421 14835 3479 14841
rect 4154 14832 4160 14844
rect 4212 14832 4218 14884
rect 4522 14832 4528 14884
rect 4580 14872 4586 14884
rect 5552 14872 5580 14903
rect 7834 14900 7840 14912
rect 7892 14900 7898 14952
rect 8202 14940 8208 14952
rect 8163 14912 8208 14940
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 11882 14900 11888 14952
rect 11940 14940 11946 14952
rect 12253 14943 12311 14949
rect 12253 14940 12265 14943
rect 11940 14912 12265 14940
rect 11940 14900 11946 14912
rect 12253 14909 12265 14912
rect 12299 14909 12311 14943
rect 13078 14940 13084 14952
rect 13039 14912 13084 14940
rect 12253 14903 12311 14909
rect 13078 14900 13084 14912
rect 13136 14900 13142 14952
rect 13446 14940 13452 14952
rect 13407 14912 13452 14940
rect 13446 14900 13452 14912
rect 13504 14900 13510 14952
rect 13725 14943 13783 14949
rect 13725 14909 13737 14943
rect 13771 14940 13783 14943
rect 14185 14943 14243 14949
rect 14185 14940 14197 14943
rect 13771 14912 14197 14940
rect 13771 14909 13783 14912
rect 13725 14903 13783 14909
rect 14185 14909 14197 14912
rect 14231 14909 14243 14943
rect 14185 14903 14243 14909
rect 14369 14943 14427 14949
rect 14369 14909 14381 14943
rect 14415 14909 14427 14943
rect 15470 14940 15476 14952
rect 15431 14912 15476 14940
rect 14369 14903 14427 14909
rect 4580 14844 5580 14872
rect 4580 14832 4586 14844
rect 9766 14832 9772 14884
rect 9824 14832 9830 14884
rect 14384 14872 14412 14903
rect 15470 14900 15476 14912
rect 15528 14900 15534 14952
rect 15749 14943 15807 14949
rect 15749 14909 15761 14943
rect 15795 14940 15807 14943
rect 16206 14940 16212 14952
rect 15795 14912 16212 14940
rect 15795 14909 15807 14912
rect 15749 14903 15807 14909
rect 16206 14900 16212 14912
rect 16264 14900 16270 14952
rect 17310 14940 17316 14952
rect 17271 14912 17316 14940
rect 17310 14900 17316 14912
rect 17368 14900 17374 14952
rect 20438 14900 20444 14952
rect 20496 14940 20502 14952
rect 20625 14943 20683 14949
rect 20625 14940 20637 14943
rect 20496 14912 20637 14940
rect 20496 14900 20502 14912
rect 20625 14909 20637 14912
rect 20671 14909 20683 14943
rect 20625 14903 20683 14909
rect 21545 14943 21603 14949
rect 21545 14909 21557 14943
rect 21591 14940 21603 14943
rect 21726 14940 21732 14952
rect 21591 14912 21732 14940
rect 21591 14909 21603 14912
rect 21545 14903 21603 14909
rect 21726 14900 21732 14912
rect 21784 14900 21790 14952
rect 24480 14943 24538 14949
rect 24480 14909 24492 14943
rect 24526 14940 24538 14943
rect 25314 14940 25320 14952
rect 24526 14912 25320 14940
rect 24526 14909 24538 14912
rect 24480 14903 24538 14909
rect 25314 14900 25320 14912
rect 25372 14900 25378 14952
rect 26510 14940 26516 14952
rect 26471 14912 26516 14940
rect 26510 14900 26516 14912
rect 26568 14900 26574 14952
rect 30926 14900 30932 14952
rect 30984 14940 30990 14952
rect 31205 14943 31263 14949
rect 31205 14940 31217 14943
rect 30984 14912 31217 14940
rect 30984 14900 30990 14912
rect 31205 14909 31217 14912
rect 31251 14909 31263 14943
rect 31386 14940 31392 14952
rect 31299 14912 31392 14940
rect 31205 14903 31263 14909
rect 31386 14900 31392 14912
rect 31444 14940 31450 14952
rect 31570 14940 31576 14952
rect 31444 14912 31576 14940
rect 31444 14900 31450 14912
rect 31570 14900 31576 14912
rect 31628 14900 31634 14952
rect 32122 14940 32128 14952
rect 32083 14912 32128 14940
rect 32122 14900 32128 14912
rect 32180 14900 32186 14952
rect 15654 14872 15660 14884
rect 14384 14844 15660 14872
rect 15654 14832 15660 14844
rect 15712 14832 15718 14884
rect 15841 14875 15899 14881
rect 15841 14841 15853 14875
rect 15887 14872 15899 14875
rect 16666 14872 16672 14884
rect 15887 14844 16672 14872
rect 15887 14841 15899 14844
rect 15841 14835 15899 14841
rect 16666 14832 16672 14844
rect 16724 14872 16730 14884
rect 20714 14872 20720 14884
rect 16724 14844 17448 14872
rect 18814 14844 20720 14872
rect 16724 14832 16730 14844
rect 17420 14816 17448 14844
rect 20714 14832 20720 14844
rect 20772 14832 20778 14884
rect 29270 14872 29276 14884
rect 29231 14844 29276 14872
rect 29270 14832 29276 14844
rect 29328 14832 29334 14884
rect 30282 14832 30288 14884
rect 30340 14832 30346 14884
rect 31297 14875 31355 14881
rect 31297 14841 31309 14875
rect 31343 14872 31355 14875
rect 31754 14872 31760 14884
rect 31343 14844 31760 14872
rect 31343 14841 31355 14844
rect 31297 14835 31355 14841
rect 31754 14832 31760 14844
rect 31812 14872 31818 14884
rect 31849 14875 31907 14881
rect 31849 14872 31861 14875
rect 31812 14844 31861 14872
rect 31812 14832 31818 14844
rect 31849 14841 31861 14844
rect 31895 14841 31907 14875
rect 31849 14835 31907 14841
rect 5169 14807 5227 14813
rect 5169 14773 5181 14807
rect 5215 14804 5227 14807
rect 5442 14804 5448 14816
rect 5215 14776 5448 14804
rect 5215 14773 5227 14776
rect 5169 14767 5227 14773
rect 5442 14764 5448 14776
rect 5500 14764 5506 14816
rect 7282 14804 7288 14816
rect 7243 14776 7288 14804
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 9033 14807 9091 14813
rect 9033 14773 9045 14807
rect 9079 14804 9091 14807
rect 11238 14804 11244 14816
rect 9079 14776 11244 14804
rect 9079 14773 9091 14776
rect 9033 14767 9091 14773
rect 11238 14764 11244 14776
rect 11296 14764 11302 14816
rect 17402 14764 17408 14816
rect 17460 14764 17466 14816
rect 19058 14804 19064 14816
rect 19019 14776 19064 14804
rect 19058 14764 19064 14776
rect 19116 14764 19122 14816
rect 20254 14764 20260 14816
rect 20312 14804 20318 14816
rect 20901 14807 20959 14813
rect 20901 14804 20913 14807
rect 20312 14776 20913 14804
rect 20312 14764 20318 14776
rect 20901 14773 20913 14776
rect 20947 14773 20959 14807
rect 21450 14804 21456 14816
rect 21411 14776 21456 14804
rect 20901 14767 20959 14773
rect 21450 14764 21456 14776
rect 21508 14764 21514 14816
rect 32033 14807 32091 14813
rect 32033 14773 32045 14807
rect 32079 14804 32091 14807
rect 32214 14804 32220 14816
rect 32079 14776 32220 14804
rect 32079 14773 32091 14776
rect 32033 14767 32091 14773
rect 32214 14764 32220 14776
rect 32272 14764 32278 14816
rect 1104 14714 34316 14736
rect 1104 14662 12052 14714
rect 12104 14662 12116 14714
rect 12168 14662 12180 14714
rect 12232 14662 12244 14714
rect 12296 14662 23123 14714
rect 23175 14662 23187 14714
rect 23239 14662 23251 14714
rect 23303 14662 23315 14714
rect 23367 14662 34316 14714
rect 1104 14640 34316 14662
rect 3145 14603 3203 14609
rect 3145 14569 3157 14603
rect 3191 14600 3203 14603
rect 3418 14600 3424 14612
rect 3191 14572 3424 14600
rect 3191 14569 3203 14572
rect 3145 14563 3203 14569
rect 3418 14560 3424 14572
rect 3476 14560 3482 14612
rect 4062 14560 4068 14612
rect 4120 14600 4126 14612
rect 4249 14603 4307 14609
rect 4249 14600 4261 14603
rect 4120 14572 4261 14600
rect 4120 14560 4126 14572
rect 4249 14569 4261 14572
rect 4295 14569 4307 14603
rect 5166 14600 5172 14612
rect 5127 14572 5172 14600
rect 4249 14563 4307 14569
rect 5166 14560 5172 14572
rect 5224 14560 5230 14612
rect 7282 14600 7288 14612
rect 5276 14572 7288 14600
rect 3329 14535 3387 14541
rect 3329 14501 3341 14535
rect 3375 14532 3387 14535
rect 4154 14532 4160 14544
rect 3375 14504 4160 14532
rect 3375 14501 3387 14504
rect 3329 14495 3387 14501
rect 4154 14492 4160 14504
rect 4212 14492 4218 14544
rect 4412 14535 4470 14541
rect 4412 14501 4424 14535
rect 4458 14532 4470 14535
rect 4522 14532 4528 14544
rect 4458 14504 4528 14532
rect 4458 14501 4470 14504
rect 4412 14495 4470 14501
rect 3053 14467 3111 14473
rect 3053 14433 3065 14467
rect 3099 14464 3111 14467
rect 4416 14464 4444 14495
rect 4522 14492 4528 14504
rect 4580 14492 4586 14544
rect 4617 14535 4675 14541
rect 4617 14501 4629 14535
rect 4663 14532 4675 14535
rect 5276 14532 5304 14572
rect 7282 14560 7288 14572
rect 7340 14560 7346 14612
rect 7377 14603 7435 14609
rect 7377 14569 7389 14603
rect 7423 14600 7435 14603
rect 7558 14600 7564 14612
rect 7423 14572 7564 14600
rect 7423 14569 7435 14572
rect 7377 14563 7435 14569
rect 7558 14560 7564 14572
rect 7616 14560 7622 14612
rect 11149 14603 11207 14609
rect 11149 14569 11161 14603
rect 11195 14600 11207 14603
rect 12710 14600 12716 14612
rect 11195 14572 12716 14600
rect 11195 14569 11207 14572
rect 11149 14563 11207 14569
rect 12710 14560 12716 14572
rect 12768 14560 12774 14612
rect 16025 14603 16083 14609
rect 16025 14569 16037 14603
rect 16071 14600 16083 14603
rect 16574 14600 16580 14612
rect 16071 14572 16580 14600
rect 16071 14569 16083 14572
rect 16025 14563 16083 14569
rect 16574 14560 16580 14572
rect 16632 14560 16638 14612
rect 20898 14600 20904 14612
rect 19996 14572 20904 14600
rect 4663 14504 5304 14532
rect 5356 14535 5414 14541
rect 4663 14501 4675 14504
rect 4617 14495 4675 14501
rect 5356 14501 5368 14535
rect 5402 14532 5414 14535
rect 5442 14532 5448 14544
rect 5402 14504 5448 14532
rect 5402 14501 5414 14504
rect 5356 14495 5414 14501
rect 5442 14492 5448 14504
rect 5500 14492 5506 14544
rect 8294 14532 8300 14544
rect 7300 14504 8300 14532
rect 5074 14464 5080 14476
rect 3099 14436 4444 14464
rect 5035 14436 5080 14464
rect 3099 14433 3111 14436
rect 3053 14427 3111 14433
rect 5074 14424 5080 14436
rect 5132 14464 5138 14476
rect 7300 14473 7328 14504
rect 8294 14492 8300 14504
rect 8352 14492 8358 14544
rect 12437 14535 12495 14541
rect 12437 14501 12449 14535
rect 12483 14532 12495 14535
rect 12802 14532 12808 14544
rect 12483 14504 12808 14532
rect 12483 14501 12495 14504
rect 12437 14495 12495 14501
rect 12802 14492 12808 14504
rect 12860 14492 12866 14544
rect 13446 14532 13452 14544
rect 13359 14504 13452 14532
rect 7285 14467 7343 14473
rect 7285 14464 7297 14467
rect 5132 14436 7297 14464
rect 5132 14424 5138 14436
rect 7285 14433 7297 14436
rect 7331 14433 7343 14467
rect 7466 14464 7472 14476
rect 7427 14436 7472 14464
rect 7285 14427 7343 14433
rect 7466 14424 7472 14436
rect 7524 14424 7530 14476
rect 11057 14467 11115 14473
rect 11057 14433 11069 14467
rect 11103 14433 11115 14467
rect 11057 14427 11115 14433
rect 11333 14467 11391 14473
rect 11333 14433 11345 14467
rect 11379 14464 11391 14467
rect 11514 14464 11520 14476
rect 11379 14436 11520 14464
rect 11379 14433 11391 14436
rect 11333 14427 11391 14433
rect 3326 14328 3332 14340
rect 3287 14300 3332 14328
rect 3326 14288 3332 14300
rect 3384 14288 3390 14340
rect 4154 14288 4160 14340
rect 4212 14328 4218 14340
rect 5353 14331 5411 14337
rect 4212 14300 4476 14328
rect 4212 14288 4218 14300
rect 4448 14269 4476 14300
rect 5353 14297 5365 14331
rect 5399 14328 5411 14331
rect 6362 14328 6368 14340
rect 5399 14300 6368 14328
rect 5399 14297 5411 14300
rect 5353 14291 5411 14297
rect 6362 14288 6368 14300
rect 6420 14288 6426 14340
rect 4433 14263 4491 14269
rect 4433 14229 4445 14263
rect 4479 14229 4491 14263
rect 11072 14260 11100 14427
rect 11514 14424 11520 14436
rect 11572 14464 11578 14476
rect 12250 14464 12256 14476
rect 11572 14436 12256 14464
rect 11572 14424 11578 14436
rect 12250 14424 12256 14436
rect 12308 14424 12314 14476
rect 12345 14467 12403 14473
rect 12345 14433 12357 14467
rect 12391 14464 12403 14467
rect 12618 14464 12624 14476
rect 12391 14436 12624 14464
rect 12391 14433 12403 14436
rect 12345 14427 12403 14433
rect 12618 14424 12624 14436
rect 12676 14424 12682 14476
rect 13372 14473 13400 14504
rect 13446 14492 13452 14504
rect 13504 14532 13510 14544
rect 13504 14504 16620 14532
rect 13504 14492 13510 14504
rect 13357 14467 13415 14473
rect 13357 14433 13369 14467
rect 13403 14433 13415 14467
rect 13357 14427 13415 14433
rect 15197 14467 15255 14473
rect 15197 14433 15209 14467
rect 15243 14464 15255 14467
rect 15286 14464 15292 14476
rect 15243 14436 15292 14464
rect 15243 14433 15255 14436
rect 15197 14427 15255 14433
rect 15286 14424 15292 14436
rect 15344 14424 15350 14476
rect 15381 14467 15439 14473
rect 15381 14433 15393 14467
rect 15427 14464 15439 14467
rect 15746 14464 15752 14476
rect 15427 14436 15752 14464
rect 15427 14433 15439 14436
rect 15381 14427 15439 14433
rect 15746 14424 15752 14436
rect 15804 14464 15810 14476
rect 16592 14473 16620 14504
rect 18414 14492 18420 14544
rect 18472 14532 18478 14544
rect 18472 14504 19012 14532
rect 18472 14492 18478 14504
rect 18984 14476 19012 14504
rect 19996 14476 20024 14572
rect 20898 14560 20904 14572
rect 20956 14560 20962 14612
rect 21726 14600 21732 14612
rect 21687 14572 21732 14600
rect 21726 14560 21732 14572
rect 21784 14600 21790 14612
rect 22278 14600 22284 14612
rect 21784 14572 22094 14600
rect 22239 14572 22284 14600
rect 21784 14560 21790 14572
rect 20254 14532 20260 14544
rect 20215 14504 20260 14532
rect 20254 14492 20260 14504
rect 20312 14492 20318 14544
rect 20714 14492 20720 14544
rect 20772 14492 20778 14544
rect 15933 14467 15991 14473
rect 15933 14464 15945 14467
rect 15804 14436 15945 14464
rect 15804 14424 15810 14436
rect 15933 14433 15945 14436
rect 15979 14433 15991 14467
rect 15933 14427 15991 14433
rect 16577 14467 16635 14473
rect 16577 14433 16589 14467
rect 16623 14433 16635 14467
rect 16758 14464 16764 14476
rect 16719 14436 16764 14464
rect 16577 14427 16635 14433
rect 16758 14424 16764 14436
rect 16816 14424 16822 14476
rect 16945 14467 17003 14473
rect 16945 14433 16957 14467
rect 16991 14464 17003 14467
rect 17954 14464 17960 14476
rect 16991 14436 17960 14464
rect 16991 14433 17003 14436
rect 16945 14427 17003 14433
rect 17954 14424 17960 14436
rect 18012 14424 18018 14476
rect 18049 14467 18107 14473
rect 18049 14433 18061 14467
rect 18095 14464 18107 14467
rect 18690 14464 18696 14476
rect 18095 14436 18696 14464
rect 18095 14433 18107 14436
rect 18049 14427 18107 14433
rect 18690 14424 18696 14436
rect 18748 14424 18754 14476
rect 18782 14424 18788 14476
rect 18840 14464 18846 14476
rect 18840 14436 18885 14464
rect 18840 14424 18846 14436
rect 18966 14424 18972 14476
rect 19024 14464 19030 14476
rect 19978 14464 19984 14476
rect 19024 14436 19117 14464
rect 19891 14436 19984 14464
rect 19024 14424 19030 14436
rect 19978 14424 19984 14436
rect 20036 14424 20042 14476
rect 22066 14464 22094 14572
rect 22278 14560 22284 14572
rect 22336 14560 22342 14612
rect 25222 14560 25228 14612
rect 25280 14600 25286 14612
rect 25317 14603 25375 14609
rect 25317 14600 25329 14603
rect 25280 14572 25329 14600
rect 25280 14560 25286 14572
rect 25317 14569 25329 14572
rect 25363 14569 25375 14603
rect 26602 14600 26608 14612
rect 25317 14563 25375 14569
rect 25424 14572 26608 14600
rect 23014 14532 23020 14544
rect 22388 14504 23020 14532
rect 22189 14467 22247 14473
rect 22189 14464 22201 14467
rect 22066 14436 22201 14464
rect 22189 14433 22201 14436
rect 22235 14433 22247 14467
rect 22189 14427 22247 14433
rect 22278 14424 22284 14476
rect 22336 14464 22342 14476
rect 22388 14473 22416 14504
rect 23014 14492 23020 14504
rect 23072 14492 23078 14544
rect 22373 14467 22431 14473
rect 22373 14464 22385 14467
rect 22336 14436 22385 14464
rect 22336 14424 22342 14436
rect 22373 14433 22385 14436
rect 22419 14433 22431 14467
rect 23032 14464 23060 14492
rect 23661 14467 23719 14473
rect 23661 14464 23673 14467
rect 23032 14436 23673 14464
rect 22373 14427 22431 14433
rect 23661 14433 23673 14436
rect 23707 14433 23719 14467
rect 23661 14427 23719 14433
rect 23845 14467 23903 14473
rect 23845 14433 23857 14467
rect 23891 14464 23903 14467
rect 24394 14464 24400 14476
rect 23891 14436 24400 14464
rect 23891 14433 23903 14436
rect 23845 14427 23903 14433
rect 24394 14424 24400 14436
rect 24452 14424 24458 14476
rect 25317 14467 25375 14473
rect 25317 14433 25329 14467
rect 25363 14464 25375 14467
rect 25424 14464 25452 14572
rect 26602 14560 26608 14572
rect 26660 14560 26666 14612
rect 27982 14560 27988 14612
rect 28040 14600 28046 14612
rect 28077 14603 28135 14609
rect 28077 14600 28089 14603
rect 28040 14572 28089 14600
rect 28040 14560 28046 14572
rect 28077 14569 28089 14572
rect 28123 14569 28135 14603
rect 28077 14563 28135 14569
rect 29270 14560 29276 14612
rect 29328 14600 29334 14612
rect 30837 14603 30895 14609
rect 30837 14600 30849 14603
rect 29328 14572 30849 14600
rect 29328 14560 29334 14572
rect 30837 14569 30849 14572
rect 30883 14569 30895 14603
rect 30837 14563 30895 14569
rect 26142 14532 26148 14544
rect 25976 14504 26148 14532
rect 25363 14436 25452 14464
rect 25501 14467 25559 14473
rect 25363 14433 25375 14436
rect 25317 14427 25375 14433
rect 25501 14433 25513 14467
rect 25547 14464 25559 14467
rect 25774 14464 25780 14476
rect 25547 14436 25780 14464
rect 25547 14433 25559 14436
rect 25501 14427 25559 14433
rect 25774 14424 25780 14436
rect 25832 14424 25838 14476
rect 25976 14473 26004 14504
rect 26142 14492 26148 14504
rect 26200 14492 26206 14544
rect 26237 14535 26295 14541
rect 26237 14501 26249 14535
rect 26283 14532 26295 14535
rect 26942 14535 27000 14541
rect 26942 14532 26954 14535
rect 26283 14504 26954 14532
rect 26283 14501 26295 14504
rect 26237 14495 26295 14501
rect 26942 14501 26954 14504
rect 26988 14501 27000 14535
rect 32030 14532 32036 14544
rect 26942 14495 27000 14501
rect 27080 14504 32036 14532
rect 25961 14467 26019 14473
rect 25961 14433 25973 14467
rect 26007 14433 26019 14467
rect 27080 14464 27108 14504
rect 32030 14492 32036 14504
rect 32088 14492 32094 14544
rect 30742 14464 30748 14476
rect 25961 14427 26019 14433
rect 26160 14436 27108 14464
rect 30703 14436 30748 14464
rect 11606 14356 11612 14408
rect 11664 14396 11670 14408
rect 12529 14399 12587 14405
rect 12529 14396 12541 14399
rect 11664 14368 12541 14396
rect 11664 14356 11670 14368
rect 12529 14365 12541 14368
rect 12575 14365 12587 14399
rect 12529 14359 12587 14365
rect 13078 14356 13084 14408
rect 13136 14396 13142 14408
rect 13173 14399 13231 14405
rect 13173 14396 13185 14399
rect 13136 14368 13185 14396
rect 13136 14356 13142 14368
rect 13173 14365 13185 14368
rect 13219 14365 13231 14399
rect 15470 14396 15476 14408
rect 15431 14368 15476 14396
rect 13173 14359 13231 14365
rect 11517 14331 11575 14337
rect 11517 14297 11529 14331
rect 11563 14328 11575 14331
rect 13188 14328 13216 14359
rect 15470 14356 15476 14368
rect 15528 14356 15534 14408
rect 18141 14399 18199 14405
rect 18141 14365 18153 14399
rect 18187 14396 18199 14399
rect 18230 14396 18236 14408
rect 18187 14368 18236 14396
rect 18187 14365 18199 14368
rect 18141 14359 18199 14365
rect 18230 14356 18236 14368
rect 18288 14356 18294 14408
rect 18325 14399 18383 14405
rect 18325 14365 18337 14399
rect 18371 14396 18383 14399
rect 18877 14399 18935 14405
rect 18877 14396 18889 14399
rect 18371 14368 18889 14396
rect 18371 14365 18383 14368
rect 18325 14359 18383 14365
rect 18877 14365 18889 14368
rect 18923 14365 18935 14399
rect 26160 14396 26188 14436
rect 30742 14424 30748 14436
rect 30800 14424 30806 14476
rect 30929 14467 30987 14473
rect 30929 14433 30941 14467
rect 30975 14464 30987 14467
rect 31938 14464 31944 14476
rect 30975 14436 31944 14464
rect 30975 14433 30987 14436
rect 30929 14427 30987 14433
rect 31938 14424 31944 14436
rect 31996 14424 32002 14476
rect 32214 14464 32220 14476
rect 32175 14436 32220 14464
rect 32214 14424 32220 14436
rect 32272 14424 32278 14476
rect 32401 14467 32459 14473
rect 32401 14433 32413 14467
rect 32447 14464 32459 14467
rect 33226 14464 33232 14476
rect 32447 14436 33232 14464
rect 32447 14433 32459 14436
rect 32401 14427 32459 14433
rect 33226 14424 33232 14436
rect 33284 14424 33290 14476
rect 18877 14359 18935 14365
rect 20088 14368 26188 14396
rect 26237 14399 26295 14405
rect 16850 14328 16856 14340
rect 11563 14300 12434 14328
rect 13188 14300 16856 14328
rect 11563 14297 11575 14300
rect 11517 14291 11575 14297
rect 11977 14263 12035 14269
rect 11977 14260 11989 14263
rect 11072 14232 11989 14260
rect 4433 14223 4491 14229
rect 11977 14229 11989 14232
rect 12023 14229 12035 14263
rect 12406 14260 12434 14300
rect 16850 14288 16856 14300
rect 16908 14288 16914 14340
rect 19058 14288 19064 14340
rect 19116 14328 19122 14340
rect 20088 14328 20116 14368
rect 26237 14365 26249 14399
rect 26283 14396 26295 14399
rect 26602 14396 26608 14408
rect 26283 14368 26608 14396
rect 26283 14365 26295 14368
rect 26237 14359 26295 14365
rect 26602 14356 26608 14368
rect 26660 14356 26666 14408
rect 26697 14399 26755 14405
rect 26697 14365 26709 14399
rect 26743 14365 26755 14399
rect 26697 14359 26755 14365
rect 23198 14328 23204 14340
rect 19116 14300 20116 14328
rect 23159 14300 23204 14328
rect 19116 14288 19122 14300
rect 23198 14288 23204 14300
rect 23256 14288 23262 14340
rect 25866 14288 25872 14340
rect 25924 14328 25930 14340
rect 26053 14331 26111 14337
rect 26053 14328 26065 14331
rect 25924 14300 26065 14328
rect 25924 14288 25930 14300
rect 26053 14297 26065 14300
rect 26099 14297 26111 14331
rect 26712 14328 26740 14359
rect 26053 14291 26111 14297
rect 26620 14300 26740 14328
rect 12710 14260 12716 14272
rect 12406 14232 12716 14260
rect 11977 14223 12035 14229
rect 12710 14220 12716 14232
rect 12768 14220 12774 14272
rect 13538 14260 13544 14272
rect 13499 14232 13544 14260
rect 13538 14220 13544 14232
rect 13596 14220 13602 14272
rect 15010 14260 15016 14272
rect 14971 14232 15016 14260
rect 15010 14220 15016 14232
rect 15068 14220 15074 14272
rect 18230 14220 18236 14272
rect 18288 14260 18294 14272
rect 23750 14260 23756 14272
rect 18288 14232 18333 14260
rect 23711 14232 23756 14260
rect 18288 14220 18294 14232
rect 23750 14220 23756 14232
rect 23808 14220 23814 14272
rect 24946 14220 24952 14272
rect 25004 14260 25010 14272
rect 26620 14260 26648 14300
rect 27614 14260 27620 14272
rect 25004 14232 27620 14260
rect 25004 14220 25010 14232
rect 27614 14220 27620 14232
rect 27672 14220 27678 14272
rect 32309 14263 32367 14269
rect 32309 14229 32321 14263
rect 32355 14260 32367 14263
rect 33318 14260 33324 14272
rect 32355 14232 33324 14260
rect 32355 14229 32367 14232
rect 32309 14223 32367 14229
rect 33318 14220 33324 14232
rect 33376 14220 33382 14272
rect 1104 14170 34316 14192
rect 1104 14118 6517 14170
rect 6569 14118 6581 14170
rect 6633 14118 6645 14170
rect 6697 14118 6709 14170
rect 6761 14118 17588 14170
rect 17640 14118 17652 14170
rect 17704 14118 17716 14170
rect 17768 14118 17780 14170
rect 17832 14118 28658 14170
rect 28710 14118 28722 14170
rect 28774 14118 28786 14170
rect 28838 14118 28850 14170
rect 28902 14118 34316 14170
rect 1104 14096 34316 14118
rect 13170 14056 13176 14068
rect 12406 14028 13176 14056
rect 8297 13991 8355 13997
rect 8297 13957 8309 13991
rect 8343 13988 8355 13991
rect 8343 13960 9260 13988
rect 8343 13957 8355 13960
rect 8297 13951 8355 13957
rect 9232 13929 9260 13960
rect 9217 13923 9275 13929
rect 9217 13889 9229 13923
rect 9263 13889 9275 13923
rect 9217 13883 9275 13889
rect 9401 13923 9459 13929
rect 9401 13889 9413 13923
rect 9447 13920 9459 13923
rect 12406 13920 12434 14028
rect 13170 14016 13176 14028
rect 13228 14056 13234 14068
rect 13630 14056 13636 14068
rect 13228 14028 13636 14056
rect 13228 14016 13234 14028
rect 13630 14016 13636 14028
rect 13688 14016 13694 14068
rect 15286 14056 15292 14068
rect 15247 14028 15292 14056
rect 15286 14016 15292 14028
rect 15344 14016 15350 14068
rect 15654 14016 15660 14068
rect 15712 14056 15718 14068
rect 16209 14059 16267 14065
rect 16209 14056 16221 14059
rect 15712 14028 16221 14056
rect 15712 14016 15718 14028
rect 16209 14025 16221 14028
rect 16255 14025 16267 14059
rect 16209 14019 16267 14025
rect 17310 14016 17316 14068
rect 17368 14056 17374 14068
rect 19978 14056 19984 14068
rect 17368 14028 19984 14056
rect 17368 14016 17374 14028
rect 17402 13988 17408 14000
rect 15580 13960 17408 13988
rect 9447 13892 12434 13920
rect 9447 13889 9459 13892
rect 9401 13883 9459 13889
rect 12894 13880 12900 13932
rect 12952 13920 12958 13932
rect 12952 13892 14136 13920
rect 12952 13880 12958 13892
rect 5442 13852 5448 13864
rect 5403 13824 5448 13852
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 5813 13855 5871 13861
rect 5813 13821 5825 13855
rect 5859 13852 5871 13855
rect 5994 13852 6000 13864
rect 5859 13824 6000 13852
rect 5859 13821 5871 13824
rect 5813 13815 5871 13821
rect 5994 13812 6000 13824
rect 6052 13812 6058 13864
rect 7009 13855 7067 13861
rect 7009 13821 7021 13855
rect 7055 13852 7067 13855
rect 7834 13852 7840 13864
rect 7055 13824 7840 13852
rect 7055 13821 7067 13824
rect 7009 13815 7067 13821
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 7926 13812 7932 13864
rect 7984 13852 7990 13864
rect 8113 13855 8171 13861
rect 8113 13852 8125 13855
rect 7984 13824 8125 13852
rect 7984 13812 7990 13824
rect 8113 13821 8125 13824
rect 8159 13821 8171 13855
rect 8113 13815 8171 13821
rect 8297 13855 8355 13861
rect 8297 13821 8309 13855
rect 8343 13852 8355 13855
rect 11606 13852 11612 13864
rect 8343 13824 11612 13852
rect 8343 13821 8355 13824
rect 8297 13815 8355 13821
rect 11606 13812 11612 13824
rect 11664 13812 11670 13864
rect 12250 13852 12256 13864
rect 12211 13824 12256 13852
rect 12250 13812 12256 13824
rect 12308 13812 12314 13864
rect 12986 13852 12992 13864
rect 12947 13824 12992 13852
rect 12986 13812 12992 13824
rect 13044 13812 13050 13864
rect 13538 13812 13544 13864
rect 13596 13852 13602 13864
rect 14108 13861 14136 13892
rect 13909 13855 13967 13861
rect 13909 13852 13921 13855
rect 13596 13824 13921 13852
rect 13596 13812 13602 13824
rect 13909 13821 13921 13824
rect 13955 13821 13967 13855
rect 13909 13815 13967 13821
rect 14093 13855 14151 13861
rect 14093 13821 14105 13855
rect 14139 13821 14151 13855
rect 14093 13815 14151 13821
rect 15378 13812 15384 13864
rect 15436 13852 15442 13864
rect 15580 13861 15608 13960
rect 17402 13948 17408 13960
rect 17460 13948 17466 14000
rect 17972 13929 18000 14028
rect 19978 14016 19984 14028
rect 20036 14016 20042 14068
rect 20809 14059 20867 14065
rect 20809 14025 20821 14059
rect 20855 14056 20867 14059
rect 20855 14028 21680 14056
rect 20855 14025 20867 14028
rect 20809 14019 20867 14025
rect 18966 13948 18972 14000
rect 19024 13988 19030 14000
rect 19337 13991 19395 13997
rect 19337 13988 19349 13991
rect 19024 13960 19349 13988
rect 19024 13948 19030 13960
rect 19337 13957 19349 13960
rect 19383 13957 19395 13991
rect 21545 13991 21603 13997
rect 21545 13988 21557 13991
rect 19337 13951 19395 13957
rect 21008 13960 21557 13988
rect 21008 13929 21036 13960
rect 21545 13957 21557 13960
rect 21591 13957 21603 13991
rect 21652 13988 21680 14028
rect 21818 14016 21824 14068
rect 21876 14056 21882 14068
rect 25590 14056 25596 14068
rect 21876 14028 25596 14056
rect 21876 14016 21882 14028
rect 25590 14016 25596 14028
rect 25648 14016 25654 14068
rect 26602 14056 26608 14068
rect 26563 14028 26608 14056
rect 26602 14016 26608 14028
rect 26660 14016 26666 14068
rect 22462 13988 22468 14000
rect 21652 13960 22468 13988
rect 21545 13951 21603 13957
rect 22462 13948 22468 13960
rect 22520 13948 22526 14000
rect 17957 13923 18015 13929
rect 17957 13889 17969 13923
rect 18003 13889 18015 13923
rect 17957 13883 18015 13889
rect 20993 13923 21051 13929
rect 20993 13889 21005 13923
rect 21039 13889 21051 13923
rect 22278 13920 22284 13932
rect 20993 13883 21051 13889
rect 21468 13892 22284 13920
rect 15746 13861 15752 13864
rect 15473 13855 15531 13861
rect 15473 13852 15485 13855
rect 15436 13824 15485 13852
rect 15436 13812 15442 13824
rect 15473 13821 15485 13824
rect 15519 13821 15531 13855
rect 15473 13815 15531 13821
rect 15565 13855 15623 13861
rect 15565 13821 15577 13855
rect 15611 13821 15623 13855
rect 15565 13815 15623 13821
rect 15693 13855 15752 13861
rect 15693 13821 15705 13855
rect 15739 13821 15752 13855
rect 15693 13815 15752 13821
rect 15746 13812 15752 13815
rect 15804 13812 15810 13864
rect 16206 13852 16212 13864
rect 16167 13824 16212 13852
rect 16206 13812 16212 13824
rect 16264 13812 16270 13864
rect 16390 13852 16396 13864
rect 16351 13824 16396 13852
rect 16390 13812 16396 13824
rect 16448 13812 16454 13864
rect 18230 13861 18236 13864
rect 18224 13852 18236 13861
rect 18191 13824 18236 13852
rect 18224 13815 18236 13824
rect 18230 13812 18236 13815
rect 18288 13812 18294 13864
rect 20717 13855 20775 13861
rect 20717 13821 20729 13855
rect 20763 13852 20775 13855
rect 20806 13852 20812 13864
rect 20763 13824 20812 13852
rect 20763 13821 20775 13824
rect 20717 13815 20775 13821
rect 20806 13812 20812 13824
rect 20864 13812 20870 13864
rect 21468 13861 21496 13892
rect 22278 13880 22284 13892
rect 22336 13880 22342 13932
rect 24394 13920 24400 13932
rect 24355 13892 24400 13920
rect 24394 13880 24400 13892
rect 24452 13880 24458 13932
rect 21453 13855 21511 13861
rect 21453 13821 21465 13855
rect 21499 13821 21511 13855
rect 21453 13815 21511 13821
rect 21637 13855 21695 13861
rect 21637 13821 21649 13855
rect 21683 13852 21695 13855
rect 21726 13852 21732 13864
rect 21683 13824 21732 13852
rect 21683 13821 21695 13824
rect 21637 13815 21695 13821
rect 21726 13812 21732 13824
rect 21784 13812 21790 13864
rect 22649 13855 22707 13861
rect 22649 13852 22661 13855
rect 22066 13824 22661 13852
rect 5000 13728 5028 13770
rect 20898 13744 20904 13796
rect 20956 13784 20962 13796
rect 22066 13784 22094 13824
rect 22649 13821 22661 13824
rect 22695 13821 22707 13855
rect 26510 13852 26516 13864
rect 26471 13824 26516 13852
rect 22649 13815 22707 13821
rect 26510 13812 26516 13824
rect 26568 13812 26574 13864
rect 26697 13855 26755 13861
rect 26697 13821 26709 13855
rect 26743 13852 26755 13855
rect 27982 13852 27988 13864
rect 26743 13824 27988 13852
rect 26743 13821 26755 13824
rect 26697 13815 26755 13821
rect 27982 13812 27988 13824
rect 28040 13812 28046 13864
rect 31205 13855 31263 13861
rect 31205 13821 31217 13855
rect 31251 13852 31263 13855
rect 31938 13852 31944 13864
rect 31251 13824 31616 13852
rect 31899 13824 31944 13852
rect 31251 13821 31263 13824
rect 31205 13815 31263 13821
rect 22922 13784 22928 13796
rect 20956 13756 22094 13784
rect 22883 13756 22928 13784
rect 20956 13744 20962 13756
rect 22922 13744 22928 13756
rect 22980 13744 22986 13796
rect 23198 13744 23204 13796
rect 23256 13784 23262 13796
rect 25038 13784 25044 13796
rect 23256 13756 23336 13784
rect 24150 13756 25044 13784
rect 23256 13744 23262 13756
rect 4062 13725 4068 13728
rect 4019 13719 4068 13725
rect 4019 13685 4031 13719
rect 4065 13685 4068 13719
rect 4019 13679 4068 13685
rect 4062 13676 4068 13679
rect 4120 13676 4126 13728
rect 4982 13676 4988 13728
rect 5040 13716 5046 13728
rect 5350 13716 5356 13728
rect 5040 13688 5356 13716
rect 5040 13676 5046 13688
rect 5350 13676 5356 13688
rect 5408 13676 5414 13728
rect 6914 13716 6920 13728
rect 6875 13688 6920 13716
rect 6914 13676 6920 13688
rect 6972 13676 6978 13728
rect 8754 13716 8760 13728
rect 8715 13688 8760 13716
rect 8754 13676 8760 13688
rect 8812 13676 8818 13728
rect 9122 13716 9128 13728
rect 9083 13688 9128 13716
rect 9122 13676 9128 13688
rect 9180 13676 9186 13728
rect 9582 13676 9588 13728
rect 9640 13716 9646 13728
rect 12529 13719 12587 13725
rect 12529 13716 12541 13719
rect 9640 13688 12541 13716
rect 9640 13676 9646 13688
rect 12529 13685 12541 13688
rect 12575 13716 12587 13719
rect 12894 13716 12900 13728
rect 12575 13688 12900 13716
rect 12575 13685 12587 13688
rect 12529 13679 12587 13685
rect 12894 13676 12900 13688
rect 12952 13676 12958 13728
rect 13906 13676 13912 13728
rect 13964 13716 13970 13728
rect 14277 13719 14335 13725
rect 14277 13716 14289 13719
rect 13964 13688 14289 13716
rect 13964 13676 13970 13688
rect 14277 13685 14289 13688
rect 14323 13685 14335 13719
rect 14277 13679 14335 13685
rect 15378 13676 15384 13728
rect 15436 13716 15442 13728
rect 16114 13716 16120 13728
rect 15436 13688 16120 13716
rect 15436 13676 15442 13688
rect 16114 13676 16120 13688
rect 16172 13676 16178 13728
rect 20990 13716 20996 13728
rect 20951 13688 20996 13716
rect 20990 13676 20996 13688
rect 21048 13676 21054 13728
rect 22830 13676 22836 13728
rect 22888 13716 22894 13728
rect 23308 13716 23336 13756
rect 25038 13744 25044 13756
rect 25096 13744 25102 13796
rect 28534 13744 28540 13796
rect 28592 13784 28598 13796
rect 30926 13784 30932 13796
rect 28592 13756 29762 13784
rect 30887 13756 30932 13784
rect 28592 13744 28598 13756
rect 30926 13744 30932 13756
rect 30984 13744 30990 13796
rect 25958 13716 25964 13728
rect 22888 13688 25964 13716
rect 22888 13676 22894 13688
rect 25958 13676 25964 13688
rect 26016 13676 26022 13728
rect 29454 13716 29460 13728
rect 29415 13688 29460 13716
rect 29454 13676 29460 13688
rect 29512 13676 29518 13728
rect 31588 13716 31616 13824
rect 31938 13812 31944 13824
rect 31996 13812 32002 13864
rect 32214 13812 32220 13864
rect 32272 13852 32278 13864
rect 33045 13855 33103 13861
rect 33045 13852 33057 13855
rect 32272 13824 33057 13852
rect 32272 13812 32278 13824
rect 33045 13821 33057 13824
rect 33091 13821 33103 13855
rect 33226 13852 33232 13864
rect 33187 13824 33232 13852
rect 33045 13815 33103 13821
rect 33226 13812 33232 13824
rect 33284 13812 33290 13864
rect 31754 13784 31760 13796
rect 31715 13756 31760 13784
rect 31754 13744 31760 13756
rect 31812 13744 31818 13796
rect 31846 13716 31852 13728
rect 31588 13688 31852 13716
rect 31846 13676 31852 13688
rect 31904 13676 31910 13728
rect 33410 13716 33416 13728
rect 33371 13688 33416 13716
rect 33410 13676 33416 13688
rect 33468 13676 33474 13728
rect 1104 13626 34316 13648
rect 1104 13574 12052 13626
rect 12104 13574 12116 13626
rect 12168 13574 12180 13626
rect 12232 13574 12244 13626
rect 12296 13574 23123 13626
rect 23175 13574 23187 13626
rect 23239 13574 23251 13626
rect 23303 13574 23315 13626
rect 23367 13574 34316 13626
rect 1104 13552 34316 13574
rect 7745 13515 7803 13521
rect 7745 13481 7757 13515
rect 7791 13512 7803 13515
rect 7834 13512 7840 13524
rect 7791 13484 7840 13512
rect 7791 13481 7803 13484
rect 7745 13475 7803 13481
rect 7834 13472 7840 13484
rect 7892 13472 7898 13524
rect 12345 13515 12403 13521
rect 12345 13512 12357 13515
rect 10336 13484 12357 13512
rect 7006 13404 7012 13456
rect 7064 13404 7070 13456
rect 10336 13453 10364 13484
rect 12345 13481 12357 13484
rect 12391 13481 12403 13515
rect 12710 13512 12716 13524
rect 12671 13484 12716 13512
rect 12345 13475 12403 13481
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 15194 13512 15200 13524
rect 12860 13484 12905 13512
rect 14752 13484 15200 13512
rect 12860 13472 12866 13484
rect 10321 13447 10379 13453
rect 10321 13413 10333 13447
rect 10367 13413 10379 13447
rect 11546 13430 13492 13444
rect 10321 13407 10379 13413
rect 11532 13416 13492 13430
rect 2866 13376 2872 13388
rect 2827 13348 2872 13376
rect 2866 13336 2872 13348
rect 2924 13336 2930 13388
rect 8573 13379 8631 13385
rect 8573 13345 8585 13379
rect 8619 13376 8631 13379
rect 8662 13376 8668 13388
rect 8619 13348 8668 13376
rect 8619 13345 8631 13348
rect 8573 13339 8631 13345
rect 8662 13336 8668 13348
rect 8720 13336 8726 13388
rect 2958 13308 2964 13320
rect 2919 13280 2964 13308
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 3050 13268 3056 13320
rect 3108 13308 3114 13320
rect 3145 13311 3203 13317
rect 3145 13308 3157 13311
rect 3108 13280 3157 13308
rect 3108 13268 3114 13280
rect 3145 13277 3157 13280
rect 3191 13308 3203 13311
rect 4706 13308 4712 13320
rect 3191 13280 4712 13308
rect 3191 13277 3203 13280
rect 3145 13271 3203 13277
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 5994 13308 6000 13320
rect 5955 13280 6000 13308
rect 5994 13268 6000 13280
rect 6052 13268 6058 13320
rect 6273 13311 6331 13317
rect 6273 13277 6285 13311
rect 6319 13308 6331 13311
rect 6914 13308 6920 13320
rect 6319 13280 6920 13308
rect 6319 13277 6331 13280
rect 6273 13271 6331 13277
rect 6914 13268 6920 13280
rect 6972 13268 6978 13320
rect 7006 13268 7012 13320
rect 7064 13308 7070 13320
rect 8018 13308 8024 13320
rect 7064 13280 8024 13308
rect 7064 13268 7070 13280
rect 8018 13268 8024 13280
rect 8076 13268 8082 13320
rect 8297 13311 8355 13317
rect 8297 13277 8309 13311
rect 8343 13308 8355 13311
rect 9950 13308 9956 13320
rect 8343 13280 9956 13308
rect 8343 13277 8355 13280
rect 8297 13271 8355 13277
rect 9950 13268 9956 13280
rect 10008 13268 10014 13320
rect 10045 13311 10103 13317
rect 10045 13277 10057 13311
rect 10091 13308 10103 13311
rect 10778 13308 10784 13320
rect 10091 13280 10784 13308
rect 10091 13277 10103 13280
rect 10045 13271 10103 13277
rect 10778 13268 10784 13280
rect 10836 13268 10842 13320
rect 10962 13268 10968 13320
rect 11020 13308 11026 13320
rect 11532 13308 11560 13416
rect 11606 13336 11612 13388
rect 11664 13376 11670 13388
rect 11664 13348 12664 13376
rect 11664 13336 11670 13348
rect 11020 13280 11560 13308
rect 11020 13268 11026 13280
rect 8481 13243 8539 13249
rect 8481 13209 8493 13243
rect 8527 13240 8539 13243
rect 8846 13240 8852 13252
rect 8527 13212 8852 13240
rect 8527 13209 8539 13212
rect 8481 13203 8539 13209
rect 8846 13200 8852 13212
rect 8904 13200 8910 13252
rect 11793 13243 11851 13249
rect 11793 13209 11805 13243
rect 11839 13240 11851 13243
rect 12636 13240 12664 13348
rect 12894 13308 12900 13320
rect 12855 13280 12900 13308
rect 12894 13268 12900 13280
rect 12952 13268 12958 13320
rect 13464 13308 13492 13416
rect 13538 13404 13544 13456
rect 13596 13444 13602 13456
rect 13725 13447 13783 13453
rect 13725 13444 13737 13447
rect 13596 13416 13737 13444
rect 13596 13404 13602 13416
rect 13725 13413 13737 13416
rect 13771 13413 13783 13447
rect 13725 13407 13783 13413
rect 13630 13336 13636 13388
rect 13688 13376 13694 13388
rect 14752 13385 14780 13484
rect 15194 13472 15200 13484
rect 15252 13472 15258 13524
rect 20714 13472 20720 13524
rect 20772 13512 20778 13524
rect 20772 13484 20852 13512
rect 20772 13472 20778 13484
rect 15010 13444 15016 13456
rect 14971 13416 15016 13444
rect 15010 13404 15016 13416
rect 15068 13404 15074 13456
rect 15286 13404 15292 13456
rect 15344 13444 15350 13456
rect 15344 13416 15502 13444
rect 15344 13404 15350 13416
rect 16758 13404 16764 13456
rect 16816 13444 16822 13456
rect 17221 13447 17279 13453
rect 17221 13444 17233 13447
rect 16816 13416 17233 13444
rect 16816 13404 16822 13416
rect 17221 13413 17233 13416
rect 17267 13413 17279 13447
rect 20824 13430 20852 13484
rect 22922 13472 22928 13524
rect 22980 13512 22986 13524
rect 23017 13515 23075 13521
rect 23017 13512 23029 13515
rect 22980 13484 23029 13512
rect 22980 13472 22986 13484
rect 23017 13481 23029 13484
rect 23063 13481 23075 13515
rect 23017 13475 23075 13481
rect 28534 13472 28540 13524
rect 28592 13512 28598 13524
rect 31297 13515 31355 13521
rect 28592 13484 30512 13512
rect 28592 13472 28598 13484
rect 26970 13444 26976 13456
rect 26931 13416 26976 13444
rect 17221 13407 17279 13413
rect 26970 13404 26976 13416
rect 27028 13404 27034 13456
rect 28813 13447 28871 13453
rect 28813 13413 28825 13447
rect 28859 13444 28871 13447
rect 30374 13444 30380 13456
rect 28859 13416 30380 13444
rect 28859 13413 28871 13416
rect 28813 13407 28871 13413
rect 30374 13404 30380 13416
rect 30432 13404 30438 13456
rect 30484 13444 30512 13484
rect 31297 13481 31309 13515
rect 31343 13512 31355 13515
rect 32214 13512 32220 13524
rect 31343 13484 32220 13512
rect 31343 13481 31355 13484
rect 31297 13475 31355 13481
rect 32214 13472 32220 13484
rect 32272 13472 32278 13524
rect 32582 13444 32588 13456
rect 30484 13416 32588 13444
rect 32582 13404 32588 13416
rect 32640 13404 32646 13456
rect 14737 13379 14795 13385
rect 14737 13376 14749 13379
rect 13688 13348 14749 13376
rect 13688 13336 13694 13348
rect 14737 13345 14749 13348
rect 14783 13345 14795 13379
rect 14737 13339 14795 13345
rect 16298 13336 16304 13388
rect 16356 13376 16362 13388
rect 17313 13379 17371 13385
rect 17313 13376 17325 13379
rect 16356 13348 17325 13376
rect 16356 13336 16362 13348
rect 17313 13345 17325 13348
rect 17359 13345 17371 13379
rect 17313 13339 17371 13345
rect 17402 13336 17408 13388
rect 17460 13376 17466 13388
rect 17589 13379 17647 13385
rect 17589 13376 17601 13379
rect 17460 13348 17601 13376
rect 17460 13336 17466 13348
rect 17589 13345 17601 13348
rect 17635 13345 17647 13379
rect 18230 13376 18236 13388
rect 18191 13348 18236 13376
rect 17589 13339 17647 13345
rect 18230 13336 18236 13348
rect 18288 13336 18294 13388
rect 18414 13376 18420 13388
rect 18375 13348 18420 13376
rect 18414 13336 18420 13348
rect 18472 13336 18478 13388
rect 18690 13336 18696 13388
rect 18748 13376 18754 13388
rect 18785 13379 18843 13385
rect 18785 13376 18797 13379
rect 18748 13348 18797 13376
rect 18748 13336 18754 13348
rect 18785 13345 18797 13348
rect 18831 13376 18843 13379
rect 18966 13376 18972 13388
rect 18831 13348 18972 13376
rect 18831 13345 18843 13348
rect 18785 13339 18843 13345
rect 18966 13336 18972 13348
rect 19024 13336 19030 13388
rect 22738 13376 22744 13388
rect 22699 13348 22744 13376
rect 22738 13336 22744 13348
rect 22796 13336 22802 13388
rect 22830 13336 22836 13388
rect 22888 13376 22894 13388
rect 23845 13379 23903 13385
rect 22888 13348 22933 13376
rect 22888 13336 22894 13348
rect 23845 13345 23857 13379
rect 23891 13376 23903 13379
rect 26142 13376 26148 13388
rect 23891 13348 26148 13376
rect 23891 13345 23903 13348
rect 23845 13339 23903 13345
rect 26142 13336 26148 13348
rect 26200 13336 26206 13388
rect 27157 13379 27215 13385
rect 27157 13345 27169 13379
rect 27203 13376 27215 13379
rect 28166 13376 28172 13388
rect 27203 13348 28172 13376
rect 27203 13345 27215 13348
rect 27157 13339 27215 13345
rect 28166 13336 28172 13348
rect 28224 13376 28230 13388
rect 28629 13379 28687 13385
rect 28629 13376 28641 13379
rect 28224 13348 28641 13376
rect 28224 13336 28230 13348
rect 28629 13345 28641 13348
rect 28675 13345 28687 13379
rect 28629 13339 28687 13345
rect 28905 13379 28963 13385
rect 28905 13345 28917 13379
rect 28951 13376 28963 13379
rect 29546 13376 29552 13388
rect 28951 13348 29552 13376
rect 28951 13345 28963 13348
rect 28905 13339 28963 13345
rect 29546 13336 29552 13348
rect 29604 13376 29610 13388
rect 30653 13379 30711 13385
rect 30653 13376 30665 13379
rect 29604 13348 30665 13376
rect 29604 13336 29610 13348
rect 30653 13345 30665 13348
rect 30699 13345 30711 13379
rect 30653 13339 30711 13345
rect 31018 13336 31024 13388
rect 31076 13376 31082 13388
rect 31205 13379 31263 13385
rect 31205 13376 31217 13379
rect 31076 13348 31217 13376
rect 31076 13336 31082 13348
rect 31205 13345 31217 13348
rect 31251 13345 31263 13379
rect 31205 13339 31263 13345
rect 15378 13308 15384 13320
rect 13464 13280 15384 13308
rect 15378 13268 15384 13280
rect 15436 13268 15442 13320
rect 15470 13268 15476 13320
rect 15528 13308 15534 13320
rect 16022 13308 16028 13320
rect 15528 13280 16028 13308
rect 15528 13268 15534 13280
rect 16022 13268 16028 13280
rect 16080 13308 16086 13320
rect 16761 13311 16819 13317
rect 16761 13308 16773 13311
rect 16080 13280 16773 13308
rect 16080 13268 16086 13280
rect 16761 13277 16773 13280
rect 16807 13277 16819 13311
rect 16761 13271 16819 13277
rect 20073 13311 20131 13317
rect 20073 13277 20085 13311
rect 20119 13308 20131 13311
rect 20349 13311 20407 13317
rect 20119 13280 20208 13308
rect 20119 13277 20131 13280
rect 20073 13271 20131 13277
rect 13541 13243 13599 13249
rect 13541 13240 13553 13243
rect 11839 13212 12434 13240
rect 12636 13212 13553 13240
rect 11839 13209 11851 13212
rect 11793 13203 11851 13209
rect 1762 13132 1768 13184
rect 1820 13172 1826 13184
rect 2501 13175 2559 13181
rect 2501 13172 2513 13175
rect 1820 13144 2513 13172
rect 1820 13132 1826 13144
rect 2501 13141 2513 13144
rect 2547 13141 2559 13175
rect 2501 13135 2559 13141
rect 7834 13132 7840 13184
rect 7892 13172 7898 13184
rect 8389 13175 8447 13181
rect 8389 13172 8401 13175
rect 7892 13144 8401 13172
rect 7892 13132 7898 13144
rect 8389 13141 8401 13144
rect 8435 13141 8447 13175
rect 8389 13135 8447 13141
rect 11054 13132 11060 13184
rect 11112 13172 11118 13184
rect 11514 13172 11520 13184
rect 11112 13144 11520 13172
rect 11112 13132 11118 13144
rect 11514 13132 11520 13144
rect 11572 13132 11578 13184
rect 12406 13172 12434 13212
rect 13541 13209 13553 13212
rect 13587 13209 13599 13243
rect 13541 13203 13599 13209
rect 13078 13172 13084 13184
rect 12406 13144 13084 13172
rect 13078 13132 13084 13144
rect 13136 13132 13142 13184
rect 20180 13172 20208 13280
rect 20349 13277 20361 13311
rect 20395 13308 20407 13311
rect 20990 13308 20996 13320
rect 20395 13280 20996 13308
rect 20395 13277 20407 13280
rect 20349 13271 20407 13277
rect 20990 13268 20996 13280
rect 21048 13268 21054 13320
rect 23017 13311 23075 13317
rect 23017 13277 23029 13311
rect 23063 13308 23075 13311
rect 23750 13308 23756 13320
rect 23063 13280 23756 13308
rect 23063 13277 23075 13280
rect 23017 13271 23075 13277
rect 23750 13268 23756 13280
rect 23808 13268 23814 13320
rect 24118 13308 24124 13320
rect 24079 13280 24124 13308
rect 24118 13268 24124 13280
rect 24176 13268 24182 13320
rect 31846 13308 31852 13320
rect 31807 13280 31852 13308
rect 31846 13268 31852 13280
rect 31904 13268 31910 13320
rect 32122 13308 32128 13320
rect 32083 13280 32128 13308
rect 32122 13268 32128 13280
rect 32180 13268 32186 13320
rect 22462 13200 22468 13252
rect 22520 13240 22526 13252
rect 23937 13243 23995 13249
rect 23937 13240 23949 13243
rect 22520 13212 23949 13240
rect 22520 13200 22526 13212
rect 23937 13209 23949 13212
rect 23983 13209 23995 13243
rect 23937 13203 23995 13209
rect 33226 13200 33232 13252
rect 33284 13240 33290 13252
rect 33597 13243 33655 13249
rect 33597 13240 33609 13243
rect 33284 13212 33609 13240
rect 33284 13200 33290 13212
rect 33597 13209 33609 13212
rect 33643 13209 33655 13243
rect 33597 13203 33655 13209
rect 20898 13172 20904 13184
rect 20180 13144 20904 13172
rect 20898 13132 20904 13144
rect 20956 13132 20962 13184
rect 21726 13132 21732 13184
rect 21784 13172 21790 13184
rect 21821 13175 21879 13181
rect 21821 13172 21833 13175
rect 21784 13144 21833 13172
rect 21784 13132 21790 13144
rect 21821 13141 21833 13144
rect 21867 13141 21879 13175
rect 21821 13135 21879 13141
rect 24026 13132 24032 13184
rect 24084 13172 24090 13184
rect 24084 13144 24129 13172
rect 24084 13132 24090 13144
rect 28074 13132 28080 13184
rect 28132 13172 28138 13184
rect 28445 13175 28503 13181
rect 28445 13172 28457 13175
rect 28132 13144 28457 13172
rect 28132 13132 28138 13144
rect 28445 13141 28457 13144
rect 28491 13141 28503 13175
rect 28445 13135 28503 13141
rect 30466 13132 30472 13184
rect 30524 13172 30530 13184
rect 30561 13175 30619 13181
rect 30561 13172 30573 13175
rect 30524 13144 30573 13172
rect 30524 13132 30530 13144
rect 30561 13141 30573 13144
rect 30607 13141 30619 13175
rect 30561 13135 30619 13141
rect 1104 13082 34316 13104
rect 1104 13030 6517 13082
rect 6569 13030 6581 13082
rect 6633 13030 6645 13082
rect 6697 13030 6709 13082
rect 6761 13030 17588 13082
rect 17640 13030 17652 13082
rect 17704 13030 17716 13082
rect 17768 13030 17780 13082
rect 17832 13030 28658 13082
rect 28710 13030 28722 13082
rect 28774 13030 28786 13082
rect 28838 13030 28850 13082
rect 28902 13030 34316 13082
rect 1104 13008 34316 13030
rect 2958 12928 2964 12980
rect 3016 12968 3022 12980
rect 3191 12971 3249 12977
rect 3191 12968 3203 12971
rect 3016 12940 3203 12968
rect 3016 12928 3022 12940
rect 3191 12937 3203 12940
rect 3237 12937 3249 12971
rect 3191 12931 3249 12937
rect 5353 12971 5411 12977
rect 5353 12937 5365 12971
rect 5399 12968 5411 12971
rect 5442 12968 5448 12980
rect 5399 12940 5448 12968
rect 5399 12937 5411 12940
rect 5353 12931 5411 12937
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 8662 12968 8668 12980
rect 8623 12940 8668 12968
rect 8662 12928 8668 12940
rect 8720 12928 8726 12980
rect 12618 12968 12624 12980
rect 12579 12940 12624 12968
rect 12618 12928 12624 12940
rect 12676 12928 12682 12980
rect 13998 12968 14004 12980
rect 13959 12940 14004 12968
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 16298 12968 16304 12980
rect 16259 12940 16304 12968
rect 16298 12928 16304 12940
rect 16356 12928 16362 12980
rect 20898 12928 20904 12980
rect 20956 12968 20962 12980
rect 21266 12968 21272 12980
rect 20956 12940 21272 12968
rect 20956 12928 20962 12940
rect 21266 12928 21272 12940
rect 21324 12968 21330 12980
rect 21637 12971 21695 12977
rect 21637 12968 21649 12971
rect 21324 12940 21649 12968
rect 21324 12928 21330 12940
rect 21637 12937 21649 12940
rect 21683 12968 21695 12971
rect 21910 12968 21916 12980
rect 21683 12940 21916 12968
rect 21683 12937 21695 12940
rect 21637 12931 21695 12937
rect 21910 12928 21916 12940
rect 21968 12928 21974 12980
rect 25038 12968 25044 12980
rect 22066 12940 25044 12968
rect 22066 12912 22094 12940
rect 25038 12928 25044 12940
rect 25096 12928 25102 12980
rect 26050 12968 26056 12980
rect 26011 12940 26056 12968
rect 26050 12928 26056 12940
rect 26108 12928 26114 12980
rect 29546 12968 29552 12980
rect 29507 12940 29552 12968
rect 29546 12928 29552 12940
rect 29604 12928 29610 12980
rect 30285 12971 30343 12977
rect 30285 12937 30297 12971
rect 30331 12968 30343 12971
rect 30926 12968 30932 12980
rect 30331 12940 30932 12968
rect 30331 12937 30343 12940
rect 30285 12931 30343 12937
rect 30926 12928 30932 12940
rect 30984 12928 30990 12980
rect 32122 12928 32128 12980
rect 32180 12968 32186 12980
rect 33045 12971 33103 12977
rect 33045 12968 33057 12971
rect 32180 12940 33057 12968
rect 32180 12928 32186 12940
rect 33045 12937 33057 12940
rect 33091 12937 33103 12971
rect 33045 12931 33103 12937
rect 9582 12900 9588 12912
rect 8128 12872 9588 12900
rect 1762 12832 1768 12844
rect 1723 12804 1768 12832
rect 1762 12792 1768 12804
rect 1820 12792 1826 12844
rect 4706 12832 4712 12844
rect 4667 12804 4712 12832
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 7926 12832 7932 12844
rect 7887 12804 7932 12832
rect 7926 12792 7932 12804
rect 7984 12792 7990 12844
rect 8128 12841 8156 12872
rect 9582 12860 9588 12872
rect 9640 12860 9646 12912
rect 10778 12860 10784 12912
rect 10836 12900 10842 12912
rect 12345 12903 12403 12909
rect 12345 12900 12357 12903
rect 10836 12872 12357 12900
rect 10836 12860 10842 12872
rect 12345 12869 12357 12872
rect 12391 12869 12403 12903
rect 13630 12900 13636 12912
rect 12345 12863 12403 12869
rect 12820 12872 13636 12900
rect 8113 12835 8171 12841
rect 8113 12801 8125 12835
rect 8159 12801 8171 12835
rect 9122 12832 9128 12844
rect 9083 12804 9128 12832
rect 8113 12795 8171 12801
rect 9122 12792 9128 12804
rect 9180 12792 9186 12844
rect 9309 12835 9367 12841
rect 9309 12801 9321 12835
rect 9355 12832 9367 12835
rect 11054 12832 11060 12844
rect 9355 12804 11060 12832
rect 9355 12801 9367 12804
rect 9309 12795 9367 12801
rect 11054 12792 11060 12804
rect 11112 12792 11118 12844
rect 12360 12832 12388 12863
rect 12820 12832 12848 12872
rect 13630 12860 13636 12872
rect 13688 12860 13694 12912
rect 18782 12900 18788 12912
rect 14108 12872 18788 12900
rect 12360 12804 12848 12832
rect 12894 12792 12900 12844
rect 12952 12832 12958 12844
rect 13170 12832 13176 12844
rect 12952 12804 13176 12832
rect 12952 12792 12958 12804
rect 13170 12792 13176 12804
rect 13228 12792 13234 12844
rect 13814 12832 13820 12844
rect 13775 12804 13820 12832
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 1394 12764 1400 12776
rect 1355 12736 1400 12764
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 4062 12724 4068 12776
rect 4120 12764 4126 12776
rect 4893 12767 4951 12773
rect 4893 12764 4905 12767
rect 4120 12736 4905 12764
rect 4120 12724 4126 12736
rect 4893 12733 4905 12736
rect 4939 12733 4951 12767
rect 7834 12764 7840 12776
rect 7795 12736 7840 12764
rect 4893 12727 4951 12733
rect 7834 12724 7840 12736
rect 7892 12724 7898 12776
rect 8754 12724 8760 12776
rect 8812 12764 8818 12776
rect 9033 12767 9091 12773
rect 9033 12764 9045 12767
rect 8812 12736 9045 12764
rect 8812 12724 8818 12736
rect 9033 12733 9045 12736
rect 9079 12733 9091 12767
rect 9033 12727 9091 12733
rect 10045 12767 10103 12773
rect 10045 12733 10057 12767
rect 10091 12764 10103 12767
rect 12161 12767 12219 12773
rect 12161 12764 12173 12767
rect 10091 12736 12173 12764
rect 10091 12733 10103 12736
rect 10045 12727 10103 12733
rect 12161 12733 12173 12736
rect 12207 12764 12219 12767
rect 12342 12764 12348 12776
rect 12207 12736 12348 12764
rect 12207 12733 12219 12736
rect 12161 12727 12219 12733
rect 12342 12724 12348 12736
rect 12400 12724 12406 12776
rect 12802 12724 12808 12776
rect 12860 12764 12866 12776
rect 12989 12767 13047 12773
rect 12989 12764 13001 12767
rect 12860 12736 13001 12764
rect 12860 12724 12866 12736
rect 12989 12733 13001 12736
rect 13035 12733 13047 12767
rect 12989 12727 13047 12733
rect 13081 12767 13139 12773
rect 13081 12733 13093 12767
rect 13127 12764 13139 12767
rect 13906 12764 13912 12776
rect 13127 12736 13912 12764
rect 13127 12733 13139 12736
rect 13081 12727 13139 12733
rect 13906 12724 13912 12736
rect 13964 12724 13970 12776
rect 14108 12773 14136 12872
rect 18782 12860 18788 12872
rect 18840 12900 18846 12912
rect 19978 12900 19984 12912
rect 18840 12872 19984 12900
rect 18840 12860 18846 12872
rect 19978 12860 19984 12872
rect 20036 12860 20042 12912
rect 20714 12860 20720 12912
rect 20772 12900 20778 12912
rect 22002 12900 22008 12912
rect 20772 12872 22008 12900
rect 20772 12860 20778 12872
rect 22002 12860 22008 12872
rect 22060 12872 22094 12912
rect 22060 12860 22066 12872
rect 22462 12860 22468 12912
rect 22520 12900 22526 12912
rect 22741 12903 22799 12909
rect 22741 12900 22753 12903
rect 22520 12872 22753 12900
rect 22520 12860 22526 12872
rect 22741 12869 22753 12872
rect 22787 12869 22799 12903
rect 26142 12900 26148 12912
rect 26103 12872 26148 12900
rect 22741 12863 22799 12869
rect 26142 12860 26148 12872
rect 26200 12860 26206 12912
rect 17954 12792 17960 12844
rect 18012 12832 18018 12844
rect 18693 12835 18751 12841
rect 18693 12832 18705 12835
rect 18012 12804 18705 12832
rect 18012 12792 18018 12804
rect 18693 12801 18705 12804
rect 18739 12801 18751 12835
rect 18693 12795 18751 12801
rect 22557 12835 22615 12841
rect 22557 12801 22569 12835
rect 22603 12832 22615 12835
rect 23566 12832 23572 12844
rect 22603 12804 23572 12832
rect 22603 12801 22615 12804
rect 22557 12795 22615 12801
rect 23566 12792 23572 12804
rect 23624 12792 23630 12844
rect 24026 12832 24032 12844
rect 23987 12804 24032 12832
rect 24026 12792 24032 12804
rect 24084 12792 24090 12844
rect 26234 12832 26240 12844
rect 26195 12804 26240 12832
rect 26234 12792 26240 12804
rect 26292 12792 26298 12844
rect 27614 12792 27620 12844
rect 27672 12832 27678 12844
rect 27798 12832 27804 12844
rect 27672 12804 27804 12832
rect 27672 12792 27678 12804
rect 27798 12792 27804 12804
rect 27856 12792 27862 12844
rect 28074 12832 28080 12844
rect 28035 12804 28080 12832
rect 28074 12792 28080 12804
rect 28132 12792 28138 12844
rect 29564 12832 29592 12928
rect 30374 12900 30380 12912
rect 30335 12872 30380 12900
rect 30374 12860 30380 12872
rect 30432 12860 30438 12912
rect 29564 12804 30972 12832
rect 14093 12767 14151 12773
rect 14093 12733 14105 12767
rect 14139 12733 14151 12767
rect 16206 12764 16212 12776
rect 16167 12736 16212 12764
rect 14093 12727 14151 12733
rect 16206 12724 16212 12736
rect 16264 12724 16270 12776
rect 16393 12767 16451 12773
rect 16393 12733 16405 12767
rect 16439 12733 16451 12767
rect 17678 12764 17684 12776
rect 17639 12736 17684 12764
rect 16393 12727 16451 12733
rect 5350 12696 5356 12708
rect 2806 12682 5356 12696
rect 2792 12668 5356 12682
rect 2682 12588 2688 12640
rect 2740 12628 2746 12640
rect 2792 12628 2820 12668
rect 5350 12656 5356 12668
rect 5408 12656 5414 12708
rect 5994 12656 6000 12708
rect 6052 12696 6058 12708
rect 6052 12668 9904 12696
rect 6052 12656 6058 12668
rect 2740 12600 2820 12628
rect 4985 12631 5043 12637
rect 2740 12588 2746 12600
rect 4985 12597 4997 12631
rect 5031 12628 5043 12631
rect 5442 12628 5448 12640
rect 5031 12600 5448 12628
rect 5031 12597 5043 12600
rect 4985 12591 5043 12597
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 7098 12588 7104 12640
rect 7156 12628 7162 12640
rect 9876 12637 9904 12668
rect 7469 12631 7527 12637
rect 7469 12628 7481 12631
rect 7156 12600 7481 12628
rect 7156 12588 7162 12600
rect 7469 12597 7481 12600
rect 7515 12597 7527 12631
rect 7469 12591 7527 12597
rect 9861 12631 9919 12637
rect 9861 12597 9873 12631
rect 9907 12597 9919 12631
rect 9861 12591 9919 12597
rect 13817 12631 13875 12637
rect 13817 12597 13829 12631
rect 13863 12628 13875 12631
rect 14642 12628 14648 12640
rect 13863 12600 14648 12628
rect 13863 12597 13875 12600
rect 13817 12591 13875 12597
rect 14642 12588 14648 12600
rect 14700 12588 14706 12640
rect 16224 12628 16252 12724
rect 16408 12696 16436 12727
rect 17678 12724 17684 12736
rect 17736 12724 17742 12776
rect 18046 12764 18052 12776
rect 18007 12736 18052 12764
rect 18046 12724 18052 12736
rect 18104 12724 18110 12776
rect 18506 12764 18512 12776
rect 18467 12736 18512 12764
rect 18506 12724 18512 12736
rect 18564 12724 18570 12776
rect 18785 12767 18843 12773
rect 18785 12733 18797 12767
rect 18831 12733 18843 12767
rect 19153 12767 19211 12773
rect 19153 12764 19165 12767
rect 18785 12727 18843 12733
rect 18892 12736 19165 12764
rect 17954 12696 17960 12708
rect 16408 12668 17960 12696
rect 17954 12656 17960 12668
rect 18012 12696 18018 12708
rect 18800 12696 18828 12727
rect 18012 12668 18828 12696
rect 18012 12656 18018 12668
rect 18892 12628 18920 12736
rect 19153 12733 19165 12736
rect 19199 12733 19211 12767
rect 19153 12727 19211 12733
rect 21821 12767 21879 12773
rect 21821 12733 21833 12767
rect 21867 12764 21879 12767
rect 22646 12764 22652 12776
rect 21867 12736 22652 12764
rect 21867 12733 21879 12736
rect 21821 12727 21879 12733
rect 22646 12724 22652 12736
rect 22704 12724 22710 12776
rect 22833 12767 22891 12773
rect 22833 12733 22845 12767
rect 22879 12733 22891 12767
rect 22833 12727 22891 12733
rect 22370 12656 22376 12708
rect 22428 12696 22434 12708
rect 22848 12696 22876 12727
rect 23014 12724 23020 12776
rect 23072 12764 23078 12776
rect 23753 12767 23811 12773
rect 23753 12764 23765 12767
rect 23072 12736 23765 12764
rect 23072 12724 23078 12736
rect 23753 12733 23765 12736
rect 23799 12733 23811 12767
rect 25958 12764 25964 12776
rect 25919 12736 25964 12764
rect 23753 12727 23811 12733
rect 25958 12724 25964 12736
rect 26016 12724 26022 12776
rect 29546 12724 29552 12776
rect 29604 12764 29610 12776
rect 30101 12767 30159 12773
rect 30101 12764 30113 12767
rect 29604 12736 30113 12764
rect 29604 12724 29610 12736
rect 30101 12733 30113 12736
rect 30147 12733 30159 12767
rect 30101 12727 30159 12733
rect 30193 12767 30251 12773
rect 30193 12733 30205 12767
rect 30239 12733 30251 12767
rect 30193 12727 30251 12733
rect 22428 12668 22876 12696
rect 22428 12656 22434 12668
rect 25038 12656 25044 12708
rect 25096 12656 25102 12708
rect 28534 12656 28540 12708
rect 28592 12656 28598 12708
rect 30208 12696 30236 12727
rect 30466 12724 30472 12776
rect 30524 12764 30530 12776
rect 30944 12773 30972 12804
rect 30929 12767 30987 12773
rect 30524 12736 30569 12764
rect 30524 12724 30530 12736
rect 30929 12733 30941 12767
rect 30975 12733 30987 12767
rect 31110 12764 31116 12776
rect 31071 12736 31116 12764
rect 30929 12727 30987 12733
rect 31110 12724 31116 12736
rect 31168 12724 31174 12776
rect 31754 12724 31760 12776
rect 31812 12764 31818 12776
rect 33045 12767 33103 12773
rect 33045 12764 33057 12767
rect 31812 12736 33057 12764
rect 31812 12724 31818 12736
rect 33045 12733 33057 12736
rect 33091 12733 33103 12767
rect 33318 12764 33324 12776
rect 33279 12736 33324 12764
rect 33045 12727 33103 12733
rect 33318 12724 33324 12736
rect 33376 12724 33382 12776
rect 30282 12696 30288 12708
rect 30195 12668 30288 12696
rect 30282 12656 30288 12668
rect 30340 12696 30346 12708
rect 30650 12696 30656 12708
rect 30340 12668 30656 12696
rect 30340 12656 30346 12668
rect 30650 12656 30656 12668
rect 30708 12656 30714 12708
rect 31294 12696 31300 12708
rect 31255 12668 31300 12696
rect 31294 12656 31300 12668
rect 31352 12656 31358 12708
rect 33229 12699 33287 12705
rect 33229 12665 33241 12699
rect 33275 12696 33287 12699
rect 33410 12696 33416 12708
rect 33275 12668 33416 12696
rect 33275 12665 33287 12668
rect 33229 12659 33287 12665
rect 33410 12656 33416 12668
rect 33468 12656 33474 12708
rect 16224 12600 18920 12628
rect 22557 12631 22615 12637
rect 22557 12597 22569 12631
rect 22603 12628 22615 12631
rect 22738 12628 22744 12640
rect 22603 12600 22744 12628
rect 22603 12597 22615 12600
rect 22557 12591 22615 12597
rect 22738 12588 22744 12600
rect 22796 12588 22802 12640
rect 24854 12588 24860 12640
rect 24912 12628 24918 12640
rect 25501 12631 25559 12637
rect 25501 12628 25513 12631
rect 24912 12600 25513 12628
rect 24912 12588 24918 12600
rect 25501 12597 25513 12600
rect 25547 12597 25559 12631
rect 25501 12591 25559 12597
rect 1104 12538 34316 12560
rect 1104 12486 12052 12538
rect 12104 12486 12116 12538
rect 12168 12486 12180 12538
rect 12232 12486 12244 12538
rect 12296 12486 23123 12538
rect 23175 12486 23187 12538
rect 23239 12486 23251 12538
rect 23303 12486 23315 12538
rect 23367 12486 34316 12538
rect 1104 12464 34316 12486
rect 2777 12427 2835 12433
rect 2777 12393 2789 12427
rect 2823 12424 2835 12427
rect 2866 12424 2872 12436
rect 2823 12396 2872 12424
rect 2823 12393 2835 12396
rect 2777 12387 2835 12393
rect 2866 12384 2872 12396
rect 2924 12384 2930 12436
rect 7926 12384 7932 12436
rect 7984 12424 7990 12436
rect 9493 12427 9551 12433
rect 9493 12424 9505 12427
rect 7984 12396 9505 12424
rect 7984 12384 7990 12396
rect 9493 12393 9505 12396
rect 9539 12393 9551 12427
rect 17678 12424 17684 12436
rect 17639 12396 17684 12424
rect 9493 12387 9551 12393
rect 17678 12384 17684 12396
rect 17736 12384 17742 12436
rect 17954 12384 17960 12436
rect 18012 12424 18018 12436
rect 18230 12424 18236 12436
rect 18012 12396 18236 12424
rect 18012 12384 18018 12396
rect 18230 12384 18236 12396
rect 18288 12384 18294 12436
rect 21910 12384 21916 12436
rect 21968 12424 21974 12436
rect 23014 12424 23020 12436
rect 21968 12396 23020 12424
rect 21968 12384 21974 12396
rect 23014 12384 23020 12396
rect 23072 12384 23078 12436
rect 23566 12424 23572 12436
rect 23527 12396 23572 12424
rect 23566 12384 23572 12396
rect 23624 12384 23630 12436
rect 24118 12424 24124 12436
rect 24079 12396 24124 12424
rect 24118 12384 24124 12396
rect 24176 12384 24182 12436
rect 25958 12424 25964 12436
rect 24228 12396 25964 12424
rect 1762 12356 1768 12368
rect 1723 12328 1768 12356
rect 1762 12316 1768 12328
rect 1820 12316 1826 12368
rect 1949 12359 2007 12365
rect 1949 12325 1961 12359
rect 1995 12356 2007 12359
rect 3878 12356 3884 12368
rect 1995 12328 3884 12356
rect 1995 12325 2007 12328
rect 1949 12319 2007 12325
rect 3878 12316 3884 12328
rect 3936 12316 3942 12368
rect 5350 12316 5356 12368
rect 5408 12316 5414 12368
rect 16853 12359 16911 12365
rect 16853 12325 16865 12359
rect 16899 12356 16911 12359
rect 18138 12356 18144 12368
rect 16899 12328 18144 12356
rect 16899 12325 16911 12328
rect 16853 12319 16911 12325
rect 18138 12316 18144 12328
rect 18196 12316 18202 12368
rect 18874 12356 18880 12368
rect 18708 12328 18880 12356
rect 3145 12291 3203 12297
rect 3145 12257 3157 12291
rect 3191 12288 3203 12291
rect 4062 12288 4068 12300
rect 3191 12260 4068 12288
rect 3191 12257 3203 12260
rect 3145 12251 3203 12257
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 8573 12291 8631 12297
rect 4632 12260 5120 12288
rect 2958 12180 2964 12232
rect 3016 12220 3022 12232
rect 3053 12223 3111 12229
rect 3053 12220 3065 12223
rect 3016 12192 3065 12220
rect 3016 12180 3022 12192
rect 3053 12189 3065 12192
rect 3099 12220 3111 12223
rect 3234 12220 3240 12232
rect 3099 12192 3240 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 3234 12180 3240 12192
rect 3292 12180 3298 12232
rect 3970 12180 3976 12232
rect 4028 12220 4034 12232
rect 4632 12229 4660 12260
rect 4617 12223 4675 12229
rect 4617 12220 4629 12223
rect 4028 12192 4629 12220
rect 4028 12180 4034 12192
rect 4617 12189 4629 12192
rect 4663 12189 4675 12223
rect 4982 12220 4988 12232
rect 4943 12192 4988 12220
rect 4617 12183 4675 12189
rect 4982 12180 4988 12192
rect 5040 12180 5046 12232
rect 5092 12220 5120 12260
rect 8573 12257 8585 12291
rect 8619 12288 8631 12291
rect 9858 12288 9864 12300
rect 8619 12260 9864 12288
rect 8619 12257 8631 12260
rect 8573 12251 8631 12257
rect 9858 12248 9864 12260
rect 9916 12248 9922 12300
rect 13078 12288 13084 12300
rect 13039 12260 13084 12288
rect 13078 12248 13084 12260
rect 13136 12248 13142 12300
rect 13265 12291 13323 12297
rect 13265 12257 13277 12291
rect 13311 12288 13323 12291
rect 13446 12288 13452 12300
rect 13311 12260 13452 12288
rect 13311 12257 13323 12260
rect 13265 12251 13323 12257
rect 13446 12248 13452 12260
rect 13504 12248 13510 12300
rect 15381 12291 15439 12297
rect 15381 12257 15393 12291
rect 15427 12288 15439 12291
rect 16758 12288 16764 12300
rect 15427 12260 16764 12288
rect 15427 12257 15439 12260
rect 15381 12251 15439 12257
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 16945 12291 17003 12297
rect 16945 12257 16957 12291
rect 16991 12257 17003 12291
rect 16945 12251 17003 12257
rect 5994 12220 6000 12232
rect 5092 12192 6000 12220
rect 5994 12180 6000 12192
rect 6052 12180 6058 12232
rect 9950 12220 9956 12232
rect 9911 12192 9956 12220
rect 9950 12180 9956 12192
rect 10008 12180 10014 12232
rect 10042 12180 10048 12232
rect 10100 12220 10106 12232
rect 15657 12223 15715 12229
rect 10100 12192 10145 12220
rect 10100 12180 10106 12192
rect 15657 12189 15669 12223
rect 15703 12220 15715 12223
rect 15746 12220 15752 12232
rect 15703 12192 15752 12220
rect 15703 12189 15715 12192
rect 15657 12183 15715 12189
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 16960 12152 16988 12251
rect 17310 12248 17316 12300
rect 17368 12288 17374 12300
rect 17589 12291 17647 12297
rect 17589 12288 17601 12291
rect 17368 12260 17601 12288
rect 17368 12248 17374 12260
rect 17589 12257 17601 12260
rect 17635 12257 17647 12291
rect 17589 12251 17647 12257
rect 17773 12291 17831 12297
rect 17773 12257 17785 12291
rect 17819 12288 17831 12291
rect 17954 12288 17960 12300
rect 17819 12260 17960 12288
rect 17819 12257 17831 12260
rect 17773 12251 17831 12257
rect 17604 12220 17632 12251
rect 17954 12248 17960 12260
rect 18012 12288 18018 12300
rect 18708 12288 18736 12328
rect 18874 12316 18880 12328
rect 18932 12316 18938 12368
rect 20070 12356 20076 12368
rect 19996 12328 20076 12356
rect 19996 12297 20024 12328
rect 20070 12316 20076 12328
rect 20128 12316 20134 12368
rect 22002 12316 22008 12368
rect 22060 12316 22066 12368
rect 22738 12356 22744 12368
rect 22699 12328 22744 12356
rect 22738 12316 22744 12328
rect 22796 12316 22802 12368
rect 18012 12260 18736 12288
rect 18785 12291 18843 12297
rect 18012 12248 18018 12260
rect 18785 12257 18797 12291
rect 18831 12257 18843 12291
rect 18785 12251 18843 12257
rect 19981 12291 20039 12297
rect 19981 12257 19993 12291
rect 20027 12257 20039 12291
rect 20162 12288 20168 12300
rect 20123 12260 20168 12288
rect 19981 12251 20039 12257
rect 18800 12220 18828 12251
rect 20162 12248 20168 12260
rect 20220 12248 20226 12300
rect 23032 12297 23060 12384
rect 23106 12316 23112 12368
rect 23164 12356 23170 12368
rect 23164 12328 23612 12356
rect 23164 12316 23170 12328
rect 23017 12291 23075 12297
rect 23017 12257 23029 12291
rect 23063 12257 23075 12291
rect 23017 12251 23075 12257
rect 23477 12291 23535 12297
rect 23477 12257 23489 12291
rect 23523 12257 23535 12291
rect 23477 12251 23535 12257
rect 17604 12192 18828 12220
rect 19061 12223 19119 12229
rect 19061 12189 19073 12223
rect 19107 12220 19119 12223
rect 20073 12223 20131 12229
rect 20073 12220 20085 12223
rect 19107 12192 20085 12220
rect 19107 12189 19119 12192
rect 19061 12183 19119 12189
rect 20073 12189 20085 12192
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 22646 12180 22652 12232
rect 22704 12220 22710 12232
rect 23106 12220 23112 12232
rect 22704 12192 23112 12220
rect 22704 12180 22710 12192
rect 23106 12180 23112 12192
rect 23164 12180 23170 12232
rect 17218 12152 17224 12164
rect 16960 12124 17224 12152
rect 17218 12112 17224 12124
rect 17276 12152 17282 12164
rect 20438 12152 20444 12164
rect 17276 12124 20444 12152
rect 17276 12112 17282 12124
rect 20438 12112 20444 12124
rect 20496 12112 20502 12164
rect 5442 12044 5448 12096
rect 5500 12084 5506 12096
rect 6411 12087 6469 12093
rect 6411 12084 6423 12087
rect 5500 12056 6423 12084
rect 5500 12044 5506 12056
rect 6411 12053 6423 12056
rect 6457 12053 6469 12087
rect 8478 12084 8484 12096
rect 8439 12056 8484 12084
rect 6411 12047 6469 12053
rect 8478 12044 8484 12056
rect 8536 12044 8542 12096
rect 13262 12084 13268 12096
rect 13223 12056 13268 12084
rect 13262 12044 13268 12056
rect 13320 12044 13326 12096
rect 15470 12084 15476 12096
rect 15431 12056 15476 12084
rect 15470 12044 15476 12056
rect 15528 12044 15534 12096
rect 15562 12044 15568 12096
rect 15620 12084 15626 12096
rect 15620 12056 15665 12084
rect 15620 12044 15626 12056
rect 18322 12044 18328 12096
rect 18380 12084 18386 12096
rect 18782 12084 18788 12096
rect 18380 12056 18788 12084
rect 18380 12044 18386 12056
rect 18782 12044 18788 12056
rect 18840 12084 18846 12096
rect 18877 12087 18935 12093
rect 18877 12084 18889 12087
rect 18840 12056 18889 12084
rect 18840 12044 18846 12056
rect 18877 12053 18889 12056
rect 18923 12053 18935 12087
rect 18877 12047 18935 12053
rect 18969 12087 19027 12093
rect 18969 12053 18981 12087
rect 19015 12084 19027 12087
rect 19058 12084 19064 12096
rect 19015 12056 19064 12084
rect 19015 12053 19027 12056
rect 18969 12047 19027 12053
rect 19058 12044 19064 12056
rect 19116 12044 19122 12096
rect 21269 12087 21327 12093
rect 21269 12053 21281 12087
rect 21315 12084 21327 12087
rect 21358 12084 21364 12096
rect 21315 12056 21364 12084
rect 21315 12053 21327 12056
rect 21269 12047 21327 12053
rect 21358 12044 21364 12056
rect 21416 12084 21422 12096
rect 23492 12084 23520 12251
rect 23584 12220 23612 12328
rect 23661 12291 23719 12297
rect 23661 12257 23673 12291
rect 23707 12288 23719 12291
rect 24121 12291 24179 12297
rect 24121 12288 24133 12291
rect 23707 12260 24133 12288
rect 23707 12257 23719 12260
rect 23661 12251 23719 12257
rect 24121 12257 24133 12260
rect 24167 12288 24179 12291
rect 24228 12288 24256 12396
rect 25958 12384 25964 12396
rect 26016 12384 26022 12436
rect 28258 12424 28264 12436
rect 27080 12396 28264 12424
rect 25869 12359 25927 12365
rect 25869 12325 25881 12359
rect 25915 12356 25927 12359
rect 26142 12356 26148 12368
rect 25915 12328 26148 12356
rect 25915 12325 25927 12328
rect 25869 12319 25927 12325
rect 26142 12316 26148 12328
rect 26200 12316 26206 12368
rect 27080 12342 27108 12396
rect 28258 12384 28264 12396
rect 28316 12424 28322 12436
rect 28534 12424 28540 12436
rect 28316 12396 28540 12424
rect 28316 12384 28322 12396
rect 28534 12384 28540 12396
rect 28592 12384 28598 12436
rect 29546 12424 29552 12436
rect 29507 12396 29552 12424
rect 29546 12384 29552 12396
rect 29604 12384 29610 12436
rect 32490 12424 32496 12436
rect 29656 12396 32496 12424
rect 29656 12356 29684 12396
rect 32490 12384 32496 12396
rect 32548 12384 32554 12436
rect 33502 12424 33508 12436
rect 33244 12396 33508 12424
rect 27172 12328 29684 12356
rect 24167 12260 24256 12288
rect 24305 12291 24363 12297
rect 24167 12257 24179 12260
rect 24121 12251 24179 12257
rect 24305 12257 24317 12291
rect 24351 12288 24363 12291
rect 24854 12288 24860 12300
rect 24351 12260 24860 12288
rect 24351 12257 24363 12260
rect 24305 12251 24363 12257
rect 24854 12248 24860 12260
rect 24912 12248 24918 12300
rect 25225 12291 25283 12297
rect 25225 12257 25237 12291
rect 25271 12257 25283 12291
rect 25225 12251 25283 12257
rect 25240 12220 25268 12251
rect 25590 12220 25596 12232
rect 23584 12192 25268 12220
rect 25551 12192 25596 12220
rect 25590 12180 25596 12192
rect 25648 12180 25654 12232
rect 25866 12180 25872 12232
rect 25924 12220 25930 12232
rect 27172 12220 27200 12328
rect 30374 12316 30380 12368
rect 30432 12356 30438 12368
rect 30469 12359 30527 12365
rect 30469 12356 30481 12359
rect 30432 12328 30481 12356
rect 30432 12316 30438 12328
rect 30469 12325 30481 12328
rect 30515 12325 30527 12359
rect 30469 12319 30527 12325
rect 32309 12359 32367 12365
rect 32309 12325 32321 12359
rect 32355 12356 32367 12359
rect 33134 12356 33140 12368
rect 32355 12328 33140 12356
rect 32355 12325 32367 12328
rect 32309 12319 32367 12325
rect 33134 12316 33140 12328
rect 33192 12316 33198 12368
rect 29365 12291 29423 12297
rect 29365 12257 29377 12291
rect 29411 12288 29423 12291
rect 29454 12288 29460 12300
rect 29411 12260 29460 12288
rect 29411 12257 29423 12260
rect 29365 12251 29423 12257
rect 29454 12248 29460 12260
rect 29512 12248 29518 12300
rect 29549 12291 29607 12297
rect 29549 12257 29561 12291
rect 29595 12288 29607 12291
rect 30282 12288 30288 12300
rect 29595 12260 30288 12288
rect 29595 12257 29607 12260
rect 29549 12251 29607 12257
rect 30282 12248 30288 12260
rect 30340 12248 30346 12300
rect 30742 12288 30748 12300
rect 30703 12260 30748 12288
rect 30742 12248 30748 12260
rect 30800 12248 30806 12300
rect 31018 12288 31024 12300
rect 30979 12260 31024 12288
rect 31018 12248 31024 12260
rect 31076 12248 31082 12300
rect 31110 12248 31116 12300
rect 31168 12288 31174 12300
rect 31168 12260 31261 12288
rect 31168 12248 31174 12260
rect 31938 12248 31944 12300
rect 31996 12288 32002 12300
rect 32125 12291 32183 12297
rect 32125 12288 32137 12291
rect 31996 12260 32137 12288
rect 31996 12248 32002 12260
rect 32125 12257 32137 12260
rect 32171 12257 32183 12291
rect 32125 12251 32183 12257
rect 32401 12291 32459 12297
rect 32401 12257 32413 12291
rect 32447 12288 32459 12291
rect 33244 12288 33272 12396
rect 33502 12384 33508 12396
rect 33560 12384 33566 12436
rect 33594 12356 33600 12368
rect 33555 12328 33600 12356
rect 33594 12316 33600 12328
rect 33652 12316 33658 12368
rect 32447 12260 33272 12288
rect 33413 12291 33471 12297
rect 32447 12257 32459 12260
rect 32401 12251 32459 12257
rect 33413 12257 33425 12291
rect 33459 12257 33471 12291
rect 33413 12251 33471 12257
rect 25924 12192 27200 12220
rect 29472 12220 29500 12248
rect 31128 12220 31156 12248
rect 29472 12192 31156 12220
rect 32140 12220 32168 12251
rect 32950 12220 32956 12232
rect 32140 12192 32956 12220
rect 25924 12180 25930 12192
rect 32950 12180 32956 12192
rect 33008 12180 33014 12232
rect 25409 12155 25467 12161
rect 25409 12121 25421 12155
rect 25455 12152 25467 12155
rect 25608 12152 25636 12180
rect 25455 12124 25636 12152
rect 25455 12121 25467 12124
rect 25409 12115 25467 12121
rect 26878 12112 26884 12164
rect 26936 12152 26942 12164
rect 33428 12152 33456 12251
rect 26936 12124 33456 12152
rect 26936 12112 26942 12124
rect 21416 12056 23520 12084
rect 21416 12044 21422 12056
rect 26602 12044 26608 12096
rect 26660 12084 26666 12096
rect 27341 12087 27399 12093
rect 27341 12084 27353 12087
rect 26660 12056 27353 12084
rect 26660 12044 26666 12056
rect 27341 12053 27353 12056
rect 27387 12053 27399 12087
rect 32122 12084 32128 12096
rect 32083 12056 32128 12084
rect 27341 12047 27399 12053
rect 32122 12044 32128 12056
rect 32180 12044 32186 12096
rect 1104 11994 34316 12016
rect 1104 11942 6517 11994
rect 6569 11942 6581 11994
rect 6633 11942 6645 11994
rect 6697 11942 6709 11994
rect 6761 11942 17588 11994
rect 17640 11942 17652 11994
rect 17704 11942 17716 11994
rect 17768 11942 17780 11994
rect 17832 11942 28658 11994
rect 28710 11942 28722 11994
rect 28774 11942 28786 11994
rect 28838 11942 28850 11994
rect 28902 11942 34316 11994
rect 1104 11920 34316 11942
rect 4982 11880 4988 11892
rect 4943 11852 4988 11880
rect 4982 11840 4988 11852
rect 5040 11840 5046 11892
rect 9122 11880 9128 11892
rect 9083 11852 9128 11880
rect 9122 11840 9128 11852
rect 9180 11840 9186 11892
rect 9858 11840 9864 11892
rect 9916 11880 9922 11892
rect 11057 11883 11115 11889
rect 11057 11880 11069 11883
rect 9916 11852 11069 11880
rect 9916 11840 9922 11852
rect 11057 11849 11069 11852
rect 11103 11849 11115 11883
rect 11057 11843 11115 11849
rect 12802 11840 12808 11892
rect 12860 11880 12866 11892
rect 12897 11883 12955 11889
rect 12897 11880 12909 11883
rect 12860 11852 12909 11880
rect 12860 11840 12866 11852
rect 12897 11849 12909 11852
rect 12943 11849 12955 11883
rect 12897 11843 12955 11849
rect 15194 11840 15200 11892
rect 15252 11880 15258 11892
rect 15252 11852 15884 11880
rect 15252 11840 15258 11852
rect 2869 11815 2927 11821
rect 2869 11781 2881 11815
rect 2915 11812 2927 11815
rect 2958 11812 2964 11824
rect 2915 11784 2964 11812
rect 2915 11781 2927 11784
rect 2869 11775 2927 11781
rect 2958 11772 2964 11784
rect 3016 11772 3022 11824
rect 8573 11815 8631 11821
rect 8573 11781 8585 11815
rect 8619 11812 8631 11815
rect 9950 11812 9956 11824
rect 8619 11784 9956 11812
rect 8619 11781 8631 11784
rect 8573 11775 8631 11781
rect 9950 11772 9956 11784
rect 10008 11772 10014 11824
rect 10042 11772 10048 11824
rect 10100 11812 10106 11824
rect 10100 11784 12434 11812
rect 10100 11772 10106 11784
rect 2685 11747 2743 11753
rect 2685 11713 2697 11747
rect 2731 11744 2743 11747
rect 3513 11747 3571 11753
rect 3513 11744 3525 11747
rect 2731 11716 3525 11744
rect 2731 11713 2743 11716
rect 2685 11707 2743 11713
rect 3513 11713 3525 11716
rect 3559 11713 3571 11747
rect 5442 11744 5448 11756
rect 5403 11716 5448 11744
rect 3513 11707 3571 11713
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 5537 11747 5595 11753
rect 5537 11713 5549 11747
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 2961 11679 3019 11685
rect 2961 11645 2973 11679
rect 3007 11676 3019 11679
rect 3050 11676 3056 11688
rect 3007 11648 3056 11676
rect 3007 11645 3019 11648
rect 2961 11639 3019 11645
rect 3050 11636 3056 11648
rect 3108 11636 3114 11688
rect 3418 11676 3424 11688
rect 3379 11648 3424 11676
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 3605 11679 3663 11685
rect 3605 11645 3617 11679
rect 3651 11645 3663 11679
rect 3605 11639 3663 11645
rect 3068 11608 3096 11636
rect 3620 11608 3648 11639
rect 5166 11636 5172 11688
rect 5224 11676 5230 11688
rect 5552 11676 5580 11707
rect 5994 11704 6000 11756
rect 6052 11744 6058 11756
rect 6825 11747 6883 11753
rect 6825 11744 6837 11747
rect 6052 11716 6837 11744
rect 6052 11704 6058 11716
rect 6825 11713 6837 11716
rect 6871 11713 6883 11747
rect 7098 11744 7104 11756
rect 7059 11716 7104 11744
rect 6825 11707 6883 11713
rect 7098 11704 7104 11716
rect 7156 11704 7162 11756
rect 9769 11747 9827 11753
rect 9769 11713 9781 11747
rect 9815 11713 9827 11747
rect 9968 11744 9996 11772
rect 12406 11744 12434 11784
rect 13541 11747 13599 11753
rect 13541 11744 13553 11747
rect 9968 11716 10548 11744
rect 12406 11716 13553 11744
rect 9769 11707 9827 11713
rect 5224 11648 5580 11676
rect 5224 11636 5230 11648
rect 8478 11636 8484 11688
rect 8536 11676 8542 11688
rect 9493 11679 9551 11685
rect 9493 11676 9505 11679
rect 8536 11648 9505 11676
rect 8536 11636 8542 11648
rect 9493 11645 9505 11648
rect 9539 11645 9551 11679
rect 9784 11676 9812 11707
rect 10042 11676 10048 11688
rect 9784 11648 10048 11676
rect 9493 11639 9551 11645
rect 10042 11636 10048 11648
rect 10100 11636 10106 11688
rect 10520 11685 10548 11716
rect 13541 11713 13553 11716
rect 13587 11744 13599 11747
rect 13630 11744 13636 11756
rect 13587 11716 13636 11744
rect 13587 11713 13599 11716
rect 13541 11707 13599 11713
rect 13630 11704 13636 11716
rect 13688 11704 13694 11756
rect 15856 11753 15884 11852
rect 16758 11840 16764 11892
rect 16816 11880 16822 11892
rect 17405 11883 17463 11889
rect 17405 11880 17417 11883
rect 16816 11852 17417 11880
rect 16816 11840 16822 11852
rect 17405 11849 17417 11852
rect 17451 11849 17463 11883
rect 17405 11843 17463 11849
rect 19242 11840 19248 11892
rect 19300 11880 19306 11892
rect 19300 11852 19932 11880
rect 19300 11840 19306 11852
rect 19904 11812 19932 11852
rect 20162 11840 20168 11892
rect 20220 11880 20226 11892
rect 20349 11883 20407 11889
rect 20349 11880 20361 11883
rect 20220 11852 20361 11880
rect 20220 11840 20226 11852
rect 20349 11849 20361 11852
rect 20395 11849 20407 11883
rect 20349 11843 20407 11849
rect 20438 11840 20444 11892
rect 20496 11880 20502 11892
rect 25866 11880 25872 11892
rect 20496 11852 25872 11880
rect 20496 11840 20502 11852
rect 25866 11840 25872 11852
rect 25924 11840 25930 11892
rect 26234 11840 26240 11892
rect 26292 11880 26298 11892
rect 26513 11883 26571 11889
rect 26513 11880 26525 11883
rect 26292 11852 26525 11880
rect 26292 11840 26298 11852
rect 26513 11849 26525 11852
rect 26559 11849 26571 11883
rect 26513 11843 26571 11849
rect 32306 11812 32312 11824
rect 19904 11784 32312 11812
rect 32306 11772 32312 11784
rect 32364 11772 32370 11824
rect 33226 11772 33232 11824
rect 33284 11772 33290 11824
rect 15841 11747 15899 11753
rect 15841 11713 15853 11747
rect 15887 11744 15899 11747
rect 16114 11744 16120 11756
rect 15887 11716 16120 11744
rect 15887 11713 15899 11716
rect 15841 11707 15899 11713
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 25590 11704 25596 11756
rect 25648 11744 25654 11756
rect 27890 11744 27896 11756
rect 25648 11716 27896 11744
rect 25648 11704 25654 11716
rect 27890 11704 27896 11716
rect 27948 11704 27954 11756
rect 31386 11744 31392 11756
rect 31347 11716 31392 11744
rect 31386 11704 31392 11716
rect 31444 11704 31450 11756
rect 33244 11744 33272 11772
rect 33152 11716 33272 11744
rect 10505 11679 10563 11685
rect 10505 11645 10517 11679
rect 10551 11676 10563 11679
rect 10686 11676 10692 11688
rect 10551 11648 10692 11676
rect 10551 11645 10563 11648
rect 10505 11639 10563 11645
rect 10686 11636 10692 11648
rect 10744 11636 10750 11688
rect 10965 11679 11023 11685
rect 10965 11645 10977 11679
rect 11011 11645 11023 11679
rect 11149 11679 11207 11685
rect 11149 11676 11161 11679
rect 10965 11639 11023 11645
rect 11072 11648 11161 11676
rect 3068 11580 3648 11608
rect 5353 11611 5411 11617
rect 5353 11577 5365 11611
rect 5399 11608 5411 11611
rect 5534 11608 5540 11620
rect 5399 11580 5540 11608
rect 5399 11577 5411 11580
rect 5353 11571 5411 11577
rect 5534 11568 5540 11580
rect 5592 11568 5598 11620
rect 8036 11552 8064 11594
rect 9766 11568 9772 11620
rect 9824 11608 9830 11620
rect 10980 11608 11008 11639
rect 9824 11580 11008 11608
rect 9824 11568 9830 11580
rect 1762 11500 1768 11552
rect 1820 11540 1826 11552
rect 2685 11543 2743 11549
rect 2685 11540 2697 11543
rect 1820 11512 2697 11540
rect 1820 11500 1826 11512
rect 2685 11509 2697 11512
rect 2731 11509 2743 11543
rect 2685 11503 2743 11509
rect 8018 11500 8024 11552
rect 8076 11500 8082 11552
rect 9585 11543 9643 11549
rect 9585 11509 9597 11543
rect 9631 11540 9643 11543
rect 9674 11540 9680 11552
rect 9631 11512 9680 11540
rect 9631 11509 9643 11512
rect 9585 11503 9643 11509
rect 9674 11500 9680 11512
rect 9732 11540 9738 11552
rect 10413 11543 10471 11549
rect 10413 11540 10425 11543
rect 9732 11512 10425 11540
rect 9732 11500 9738 11512
rect 10413 11509 10425 11512
rect 10459 11509 10471 11543
rect 10413 11503 10471 11509
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11072 11540 11100 11648
rect 11149 11645 11161 11648
rect 11195 11645 11207 11679
rect 11149 11639 11207 11645
rect 15562 11636 15568 11688
rect 15620 11685 15626 11688
rect 15620 11676 15632 11685
rect 17497 11679 17555 11685
rect 15620 11648 15665 11676
rect 15620 11639 15632 11648
rect 17497 11645 17509 11679
rect 17543 11676 17555 11679
rect 18506 11676 18512 11688
rect 17543 11648 18512 11676
rect 17543 11645 17555 11648
rect 17497 11639 17555 11645
rect 15620 11636 15626 11639
rect 18506 11636 18512 11648
rect 18564 11636 18570 11688
rect 18969 11679 19027 11685
rect 18969 11645 18981 11679
rect 19015 11645 19027 11679
rect 18969 11639 19027 11645
rect 13265 11611 13323 11617
rect 13265 11577 13277 11611
rect 13311 11608 13323 11611
rect 14366 11608 14372 11620
rect 13311 11580 14372 11608
rect 13311 11577 13323 11580
rect 13265 11571 13323 11577
rect 14366 11568 14372 11580
rect 14424 11568 14430 11620
rect 18984 11608 19012 11639
rect 19058 11636 19064 11688
rect 19116 11676 19122 11688
rect 19225 11679 19283 11685
rect 19225 11676 19237 11679
rect 19116 11648 19237 11676
rect 19116 11636 19122 11648
rect 19225 11645 19237 11648
rect 19271 11645 19283 11679
rect 19225 11639 19283 11645
rect 24397 11679 24455 11685
rect 24397 11645 24409 11679
rect 24443 11676 24455 11679
rect 24854 11676 24860 11688
rect 24443 11648 24860 11676
rect 24443 11645 24455 11648
rect 24397 11639 24455 11645
rect 24854 11636 24860 11648
rect 24912 11636 24918 11688
rect 25038 11676 25044 11688
rect 24999 11648 25044 11676
rect 25038 11636 25044 11648
rect 25096 11636 25102 11688
rect 25958 11636 25964 11688
rect 26016 11676 26022 11688
rect 26421 11679 26479 11685
rect 26421 11676 26433 11679
rect 26016 11648 26433 11676
rect 26016 11636 26022 11648
rect 26421 11645 26433 11648
rect 26467 11645 26479 11679
rect 26602 11676 26608 11688
rect 26563 11648 26608 11676
rect 26421 11639 26479 11645
rect 26602 11636 26608 11648
rect 26660 11636 26666 11688
rect 28166 11676 28172 11688
rect 28127 11648 28172 11676
rect 28166 11636 28172 11648
rect 28224 11636 28230 11688
rect 28442 11676 28448 11688
rect 28403 11648 28448 11676
rect 28442 11636 28448 11648
rect 28500 11636 28506 11688
rect 29546 11676 29552 11688
rect 29507 11648 29552 11676
rect 29546 11636 29552 11648
rect 29604 11636 29610 11688
rect 29733 11679 29791 11685
rect 29733 11645 29745 11679
rect 29779 11676 29791 11679
rect 30374 11676 30380 11688
rect 29779 11648 30380 11676
rect 29779 11645 29791 11648
rect 29733 11639 29791 11645
rect 30374 11636 30380 11648
rect 30432 11636 30438 11688
rect 30742 11676 30748 11688
rect 30703 11648 30748 11676
rect 30742 11636 30748 11648
rect 30800 11636 30806 11688
rect 31018 11636 31024 11688
rect 31076 11676 31082 11688
rect 31113 11679 31171 11685
rect 31113 11676 31125 11679
rect 31076 11648 31125 11676
rect 31076 11636 31082 11648
rect 31113 11645 31125 11648
rect 31159 11645 31171 11679
rect 31113 11639 31171 11645
rect 31294 11636 31300 11688
rect 31352 11676 31358 11688
rect 33152 11685 33180 11716
rect 31481 11679 31539 11685
rect 31481 11676 31493 11679
rect 31352 11648 31493 11676
rect 31352 11636 31358 11648
rect 31481 11645 31493 11648
rect 31527 11645 31539 11679
rect 31481 11639 31539 11645
rect 33137 11679 33195 11685
rect 33137 11645 33149 11679
rect 33183 11645 33195 11679
rect 33137 11639 33195 11645
rect 33226 11636 33232 11688
rect 33284 11676 33290 11688
rect 33321 11679 33379 11685
rect 33321 11676 33333 11679
rect 33284 11648 33333 11676
rect 33284 11636 33290 11648
rect 33321 11645 33333 11648
rect 33367 11645 33379 11679
rect 33321 11639 33379 11645
rect 21266 11608 21272 11620
rect 18984 11580 21272 11608
rect 21266 11568 21272 11580
rect 21324 11568 21330 11620
rect 25777 11611 25835 11617
rect 25777 11577 25789 11611
rect 25823 11608 25835 11611
rect 28258 11608 28264 11620
rect 25823 11580 28264 11608
rect 25823 11577 25835 11580
rect 25777 11571 25835 11577
rect 28258 11568 28264 11580
rect 28316 11568 28322 11620
rect 11790 11540 11796 11552
rect 10928 11512 11796 11540
rect 10928 11500 10934 11512
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 13078 11500 13084 11552
rect 13136 11540 13142 11552
rect 13357 11543 13415 11549
rect 13357 11540 13369 11543
rect 13136 11512 13369 11540
rect 13136 11500 13142 11512
rect 13357 11509 13369 11512
rect 13403 11540 13415 11543
rect 13722 11540 13728 11552
rect 13403 11512 13728 11540
rect 13403 11509 13415 11512
rect 13357 11503 13415 11509
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 14458 11540 14464 11552
rect 14419 11512 14464 11540
rect 14458 11500 14464 11512
rect 14516 11500 14522 11552
rect 23566 11500 23572 11552
rect 23624 11540 23630 11552
rect 24305 11543 24363 11549
rect 24305 11540 24317 11543
rect 23624 11512 24317 11540
rect 23624 11500 23630 11512
rect 24305 11509 24317 11512
rect 24351 11509 24363 11543
rect 24305 11503 24363 11509
rect 27798 11500 27804 11552
rect 27856 11540 27862 11552
rect 27985 11543 28043 11549
rect 27985 11540 27997 11543
rect 27856 11512 27997 11540
rect 27856 11500 27862 11512
rect 27985 11509 27997 11512
rect 28031 11509 28043 11543
rect 27985 11503 28043 11509
rect 28353 11543 28411 11549
rect 28353 11509 28365 11543
rect 28399 11540 28411 11543
rect 29641 11543 29699 11549
rect 29641 11540 29653 11543
rect 28399 11512 29653 11540
rect 28399 11509 28411 11512
rect 28353 11503 28411 11509
rect 29641 11509 29653 11512
rect 29687 11509 29699 11543
rect 33318 11540 33324 11552
rect 33279 11512 33324 11540
rect 29641 11503 29699 11509
rect 33318 11500 33324 11512
rect 33376 11500 33382 11552
rect 1104 11450 34316 11472
rect 1104 11398 12052 11450
rect 12104 11398 12116 11450
rect 12168 11398 12180 11450
rect 12232 11398 12244 11450
rect 12296 11398 23123 11450
rect 23175 11398 23187 11450
rect 23239 11398 23251 11450
rect 23303 11398 23315 11450
rect 23367 11398 34316 11450
rect 1104 11376 34316 11398
rect 9493 11339 9551 11345
rect 9493 11305 9505 11339
rect 9539 11336 9551 11339
rect 9766 11336 9772 11348
rect 9539 11308 9772 11336
rect 9539 11305 9551 11308
rect 9493 11299 9551 11305
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 9876 11308 12434 11336
rect 2682 11228 2688 11280
rect 2740 11228 2746 11280
rect 9674 11268 9680 11280
rect 9635 11240 9680 11268
rect 9674 11228 9680 11240
rect 9732 11228 9738 11280
rect 9876 11277 9904 11308
rect 9861 11271 9919 11277
rect 9861 11237 9873 11271
rect 9907 11237 9919 11271
rect 10778 11268 10784 11280
rect 9861 11231 9919 11237
rect 10428 11240 10784 11268
rect 1394 11200 1400 11212
rect 1355 11172 1400 11200
rect 1394 11160 1400 11172
rect 1452 11160 1458 11212
rect 1762 11200 1768 11212
rect 1723 11172 1768 11200
rect 1762 11160 1768 11172
rect 1820 11160 1826 11212
rect 5258 11200 5264 11212
rect 5219 11172 5264 11200
rect 5258 11160 5264 11172
rect 5316 11160 5322 11212
rect 5353 11203 5411 11209
rect 5353 11169 5365 11203
rect 5399 11200 5411 11203
rect 5534 11200 5540 11212
rect 5399 11172 5540 11200
rect 5399 11169 5411 11172
rect 5353 11163 5411 11169
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 10428 11209 10456 11240
rect 10778 11228 10784 11240
rect 10836 11228 10842 11280
rect 11146 11228 11152 11280
rect 11204 11228 11210 11280
rect 12406 11268 12434 11308
rect 13262 11296 13268 11348
rect 13320 11336 13326 11348
rect 14900 11339 14958 11345
rect 14900 11336 14912 11339
rect 13320 11308 14912 11336
rect 13320 11296 13326 11308
rect 14900 11305 14912 11308
rect 14946 11305 14958 11339
rect 15746 11336 15752 11348
rect 15707 11308 15752 11336
rect 14900 11299 14958 11305
rect 15746 11296 15752 11308
rect 15804 11296 15810 11348
rect 18046 11336 18052 11348
rect 18007 11308 18052 11336
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 19978 11296 19984 11348
rect 20036 11336 20042 11348
rect 20625 11339 20683 11345
rect 20625 11336 20637 11339
rect 20036 11308 20637 11336
rect 20036 11296 20042 11308
rect 20625 11305 20637 11308
rect 20671 11305 20683 11339
rect 20625 11299 20683 11305
rect 23014 11296 23020 11348
rect 23072 11336 23078 11348
rect 23201 11339 23259 11345
rect 23201 11336 23213 11339
rect 23072 11308 23213 11336
rect 23072 11296 23078 11308
rect 23201 11305 23213 11308
rect 23247 11305 23259 11339
rect 23201 11299 23259 11305
rect 30561 11339 30619 11345
rect 30561 11305 30573 11339
rect 30607 11336 30619 11339
rect 31018 11336 31024 11348
rect 30607 11308 31024 11336
rect 30607 11305 30619 11308
rect 30561 11299 30619 11305
rect 31018 11296 31024 11308
rect 31076 11296 31082 11348
rect 12406 11240 13860 11268
rect 10413 11203 10471 11209
rect 10413 11169 10425 11203
rect 10459 11169 10471 11203
rect 12713 11203 12771 11209
rect 12713 11200 12725 11203
rect 10413 11163 10471 11169
rect 11900 11172 12725 11200
rect 1412 11132 1440 11160
rect 2866 11132 2872 11144
rect 1412 11104 2872 11132
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 3050 11092 3056 11144
rect 3108 11132 3114 11144
rect 5166 11132 5172 11144
rect 3108 11104 5172 11132
rect 3108 11092 3114 11104
rect 5166 11092 5172 11104
rect 5224 11132 5230 11144
rect 5445 11135 5503 11141
rect 5445 11132 5457 11135
rect 5224 11104 5457 11132
rect 5224 11092 5230 11104
rect 5445 11101 5457 11104
rect 5491 11101 5503 11135
rect 5445 11095 5503 11101
rect 10686 11092 10692 11144
rect 10744 11132 10750 11144
rect 11900 11132 11928 11172
rect 12713 11169 12725 11172
rect 12759 11169 12771 11203
rect 12713 11163 12771 11169
rect 13446 11160 13452 11212
rect 13504 11200 13510 11212
rect 13541 11203 13599 11209
rect 13541 11200 13553 11203
rect 13504 11172 13553 11200
rect 13504 11160 13510 11172
rect 13541 11169 13553 11172
rect 13587 11169 13599 11203
rect 13722 11200 13728 11212
rect 13683 11172 13728 11200
rect 13541 11163 13599 11169
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 10744 11104 11928 11132
rect 12161 11135 12219 11141
rect 10744 11092 10750 11104
rect 12161 11101 12173 11135
rect 12207 11132 12219 11135
rect 13464 11132 13492 11160
rect 12207 11104 13492 11132
rect 12207 11101 12219 11104
rect 12161 11095 12219 11101
rect 13262 11024 13268 11076
rect 13320 11064 13326 11076
rect 13541 11067 13599 11073
rect 13541 11064 13553 11067
rect 13320 11036 13553 11064
rect 13320 11024 13326 11036
rect 13541 11033 13553 11036
rect 13587 11033 13599 11067
rect 13832 11064 13860 11240
rect 14090 11228 14096 11280
rect 14148 11268 14154 11280
rect 15105 11271 15163 11277
rect 15105 11268 15117 11271
rect 14148 11240 15117 11268
rect 14148 11228 14154 11240
rect 15105 11237 15117 11240
rect 15151 11237 15163 11271
rect 18506 11268 18512 11280
rect 15105 11231 15163 11237
rect 16960 11240 18512 11268
rect 14458 11160 14464 11212
rect 14516 11200 14522 11212
rect 15657 11203 15715 11209
rect 15657 11200 15669 11203
rect 14516 11172 15669 11200
rect 14516 11160 14522 11172
rect 15657 11169 15669 11172
rect 15703 11169 15715 11203
rect 15838 11200 15844 11212
rect 15799 11172 15844 11200
rect 15657 11163 15715 11169
rect 15838 11160 15844 11172
rect 15896 11160 15902 11212
rect 16960 11209 16988 11240
rect 18506 11228 18512 11240
rect 18564 11228 18570 11280
rect 26053 11271 26111 11277
rect 26053 11237 26065 11271
rect 26099 11268 26111 11271
rect 26878 11268 26884 11280
rect 26099 11240 26884 11268
rect 26099 11237 26111 11240
rect 26053 11231 26111 11237
rect 26878 11228 26884 11240
rect 26936 11228 26942 11280
rect 27798 11268 27804 11280
rect 27759 11240 27804 11268
rect 27798 11228 27804 11240
rect 27856 11228 27862 11280
rect 28258 11228 28264 11280
rect 28316 11228 28322 11280
rect 32122 11268 32128 11280
rect 32083 11240 32128 11268
rect 32122 11228 32128 11240
rect 32180 11228 32186 11280
rect 32582 11228 32588 11280
rect 32640 11228 32646 11280
rect 16945 11203 17003 11209
rect 16945 11169 16957 11203
rect 16991 11169 17003 11203
rect 16945 11163 17003 11169
rect 18049 11203 18107 11209
rect 18049 11169 18061 11203
rect 18095 11200 18107 11203
rect 18138 11200 18144 11212
rect 18095 11172 18144 11200
rect 18095 11169 18107 11172
rect 18049 11163 18107 11169
rect 18138 11160 18144 11172
rect 18196 11160 18202 11212
rect 18233 11203 18291 11209
rect 18233 11169 18245 11203
rect 18279 11169 18291 11203
rect 18233 11163 18291 11169
rect 19061 11203 19119 11209
rect 19061 11169 19073 11203
rect 19107 11200 19119 11203
rect 19794 11200 19800 11212
rect 19107 11172 19800 11200
rect 19107 11169 19119 11172
rect 19061 11163 19119 11169
rect 18248 11132 18276 11163
rect 19794 11160 19800 11172
rect 19852 11160 19858 11212
rect 20346 11160 20352 11212
rect 20404 11200 20410 11212
rect 20441 11203 20499 11209
rect 20441 11200 20453 11203
rect 20404 11172 20453 11200
rect 20404 11160 20410 11172
rect 20441 11169 20453 11172
rect 20487 11169 20499 11203
rect 21726 11200 21732 11212
rect 21687 11172 21732 11200
rect 20441 11163 20499 11169
rect 21726 11160 21732 11172
rect 21784 11160 21790 11212
rect 22370 11200 22376 11212
rect 22331 11172 22376 11200
rect 22370 11160 22376 11172
rect 22428 11160 22434 11212
rect 22554 11200 22560 11212
rect 22515 11172 22560 11200
rect 22554 11160 22560 11172
rect 22612 11160 22618 11212
rect 22830 11160 22836 11212
rect 22888 11200 22894 11212
rect 23017 11203 23075 11209
rect 23017 11200 23029 11203
rect 22888 11172 23029 11200
rect 22888 11160 22894 11172
rect 23017 11169 23029 11172
rect 23063 11169 23075 11203
rect 23566 11200 23572 11212
rect 23527 11172 23572 11200
rect 23017 11163 23075 11169
rect 23566 11160 23572 11172
rect 23624 11160 23630 11212
rect 25682 11160 25688 11212
rect 25740 11200 25746 11212
rect 25740 11172 26280 11200
rect 25740 11160 25746 11172
rect 19242 11132 19248 11144
rect 18248 11104 19248 11132
rect 19242 11092 19248 11104
rect 19300 11092 19306 11144
rect 23842 11132 23848 11144
rect 23803 11104 23848 11132
rect 23842 11092 23848 11104
rect 23900 11092 23906 11144
rect 25958 11092 25964 11144
rect 26016 11132 26022 11144
rect 26252 11141 26280 11172
rect 26602 11160 26608 11212
rect 26660 11200 26666 11212
rect 27065 11203 27123 11209
rect 27065 11200 27077 11203
rect 26660 11172 27077 11200
rect 26660 11160 26666 11172
rect 27065 11169 27077 11172
rect 27111 11169 27123 11203
rect 30469 11203 30527 11209
rect 30469 11200 30481 11203
rect 27065 11163 27123 11169
rect 29288 11172 30481 11200
rect 26145 11135 26203 11141
rect 26145 11132 26157 11135
rect 26016 11104 26157 11132
rect 26016 11092 26022 11104
rect 26145 11101 26157 11104
rect 26191 11101 26203 11135
rect 26145 11095 26203 11101
rect 26237 11135 26295 11141
rect 26237 11101 26249 11135
rect 26283 11101 26295 11135
rect 26237 11095 26295 11101
rect 27525 11135 27583 11141
rect 27525 11101 27537 11135
rect 27571 11132 27583 11135
rect 27890 11132 27896 11144
rect 27571 11104 27896 11132
rect 27571 11101 27583 11104
rect 27525 11095 27583 11101
rect 27890 11092 27896 11104
rect 27948 11092 27954 11144
rect 29086 11092 29092 11144
rect 29144 11132 29150 11144
rect 29288 11141 29316 11172
rect 30469 11169 30481 11172
rect 30515 11169 30527 11203
rect 30469 11163 30527 11169
rect 31202 11160 31208 11212
rect 31260 11200 31266 11212
rect 31297 11203 31355 11209
rect 31297 11200 31309 11203
rect 31260 11172 31309 11200
rect 31260 11160 31266 11172
rect 31297 11169 31309 11172
rect 31343 11169 31355 11203
rect 31846 11200 31852 11212
rect 31807 11172 31852 11200
rect 31297 11163 31355 11169
rect 31846 11160 31852 11172
rect 31904 11160 31910 11212
rect 29273 11135 29331 11141
rect 29273 11132 29285 11135
rect 29144 11104 29285 11132
rect 29144 11092 29150 11104
rect 29273 11101 29285 11104
rect 29319 11101 29331 11135
rect 29273 11095 29331 11101
rect 14182 11064 14188 11076
rect 13832 11036 14188 11064
rect 13541 11027 13599 11033
rect 14182 11024 14188 11036
rect 14240 11064 14246 11076
rect 14737 11067 14795 11073
rect 14737 11064 14749 11067
rect 14240 11036 14749 11064
rect 14240 11024 14246 11036
rect 14737 11033 14749 11036
rect 14783 11033 14795 11067
rect 14737 11027 14795 11033
rect 18414 11024 18420 11076
rect 18472 11064 18478 11076
rect 18966 11064 18972 11076
rect 18472 11036 18972 11064
rect 18472 11024 18478 11036
rect 18966 11024 18972 11036
rect 19024 11024 19030 11076
rect 21542 11024 21548 11076
rect 21600 11064 21606 11076
rect 21821 11067 21879 11073
rect 21821 11064 21833 11067
rect 21600 11036 21833 11064
rect 21600 11024 21606 11036
rect 21821 11033 21833 11036
rect 21867 11033 21879 11067
rect 21821 11027 21879 11033
rect 21910 11024 21916 11076
rect 21968 11064 21974 11076
rect 22465 11067 22523 11073
rect 22465 11064 22477 11067
rect 21968 11036 22477 11064
rect 21968 11024 21974 11036
rect 22465 11033 22477 11036
rect 22511 11033 22523 11067
rect 22465 11027 22523 11033
rect 23474 11024 23480 11076
rect 23532 11064 23538 11076
rect 23661 11067 23719 11073
rect 23661 11064 23673 11067
rect 23532 11036 23673 11064
rect 23532 11024 23538 11036
rect 23661 11033 23673 11036
rect 23707 11033 23719 11067
rect 26970 11064 26976 11076
rect 26931 11036 26976 11064
rect 23661 11027 23719 11033
rect 26970 11024 26976 11036
rect 27028 11024 27034 11076
rect 2774 10956 2780 11008
rect 2832 10996 2838 11008
rect 3191 10999 3249 11005
rect 3191 10996 3203 10999
rect 2832 10968 3203 10996
rect 2832 10956 2838 10968
rect 3191 10965 3203 10968
rect 3237 10996 3249 10999
rect 3418 10996 3424 11008
rect 3237 10968 3424 10996
rect 3237 10965 3249 10968
rect 3191 10959 3249 10965
rect 3418 10956 3424 10968
rect 3476 10956 3482 11008
rect 4890 10996 4896 11008
rect 4851 10968 4896 10996
rect 4890 10956 4896 10968
rect 4948 10956 4954 11008
rect 10410 10956 10416 11008
rect 10468 10996 10474 11008
rect 10670 10999 10728 11005
rect 10670 10996 10682 10999
rect 10468 10968 10682 10996
rect 10468 10956 10474 10968
rect 10670 10965 10682 10968
rect 10716 10965 10728 10999
rect 14918 10996 14924 11008
rect 14879 10968 14924 10996
rect 10670 10959 10728 10965
rect 14918 10956 14924 10968
rect 14976 10956 14982 11008
rect 17218 10996 17224 11008
rect 17179 10968 17224 10996
rect 17218 10956 17224 10968
rect 17276 10956 17282 11008
rect 17402 10996 17408 11008
rect 17363 10968 17408 10996
rect 17402 10956 17408 10968
rect 17460 10956 17466 11008
rect 23750 10996 23756 11008
rect 23711 10968 23756 10996
rect 23750 10956 23756 10968
rect 23808 10956 23814 11008
rect 25406 10956 25412 11008
rect 25464 10996 25470 11008
rect 25685 10999 25743 11005
rect 25685 10996 25697 10999
rect 25464 10968 25697 10996
rect 25464 10956 25470 10968
rect 25685 10965 25697 10968
rect 25731 10965 25743 10999
rect 25685 10959 25743 10965
rect 28442 10956 28448 11008
rect 28500 10996 28506 11008
rect 29638 10996 29644 11008
rect 28500 10968 29644 10996
rect 28500 10956 28506 10968
rect 29638 10956 29644 10968
rect 29696 10956 29702 11008
rect 30650 10956 30656 11008
rect 30708 10996 30714 11008
rect 31205 10999 31263 11005
rect 31205 10996 31217 10999
rect 30708 10968 31217 10996
rect 30708 10956 30714 10968
rect 31205 10965 31217 10968
rect 31251 10965 31263 10999
rect 31205 10959 31263 10965
rect 33226 10956 33232 11008
rect 33284 10996 33290 11008
rect 33597 10999 33655 11005
rect 33597 10996 33609 10999
rect 33284 10968 33609 10996
rect 33284 10956 33290 10968
rect 33597 10965 33609 10968
rect 33643 10965 33655 10999
rect 33597 10959 33655 10965
rect 1104 10906 34316 10928
rect 1104 10854 6517 10906
rect 6569 10854 6581 10906
rect 6633 10854 6645 10906
rect 6697 10854 6709 10906
rect 6761 10854 17588 10906
rect 17640 10854 17652 10906
rect 17704 10854 17716 10906
rect 17768 10854 17780 10906
rect 17832 10854 28658 10906
rect 28710 10854 28722 10906
rect 28774 10854 28786 10906
rect 28838 10854 28850 10906
rect 28902 10854 34316 10906
rect 1104 10832 34316 10854
rect 3050 10752 3056 10804
rect 3108 10792 3114 10804
rect 3329 10795 3387 10801
rect 3329 10792 3341 10795
rect 3108 10764 3341 10792
rect 3108 10752 3114 10764
rect 3329 10761 3341 10764
rect 3375 10761 3387 10795
rect 3329 10755 3387 10761
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 5767 10795 5825 10801
rect 5767 10792 5779 10795
rect 5592 10764 5779 10792
rect 5592 10752 5598 10764
rect 5767 10761 5779 10764
rect 5813 10761 5825 10795
rect 5767 10755 5825 10761
rect 9769 10795 9827 10801
rect 9769 10761 9781 10795
rect 9815 10792 9827 10795
rect 10042 10792 10048 10804
rect 9815 10764 10048 10792
rect 9815 10761 9827 10764
rect 9769 10755 9827 10761
rect 10042 10752 10048 10764
rect 10100 10752 10106 10804
rect 10410 10792 10416 10804
rect 10371 10764 10416 10792
rect 10410 10752 10416 10764
rect 10468 10752 10474 10804
rect 12069 10795 12127 10801
rect 12069 10761 12081 10795
rect 12115 10792 12127 10795
rect 12342 10792 12348 10804
rect 12115 10764 12348 10792
rect 12115 10761 12127 10764
rect 12069 10755 12127 10761
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 13354 10792 13360 10804
rect 13315 10764 13360 10792
rect 13354 10752 13360 10764
rect 13412 10752 13418 10804
rect 14366 10792 14372 10804
rect 14327 10764 14372 10792
rect 14366 10752 14372 10764
rect 14424 10752 14430 10804
rect 15289 10795 15347 10801
rect 15289 10761 15301 10795
rect 15335 10792 15347 10795
rect 15470 10792 15476 10804
rect 15335 10764 15476 10792
rect 15335 10761 15347 10764
rect 15289 10755 15347 10761
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 16390 10752 16396 10804
rect 16448 10792 16454 10804
rect 18322 10792 18328 10804
rect 16448 10764 18328 10792
rect 16448 10752 16454 10764
rect 18322 10752 18328 10764
rect 18380 10752 18386 10804
rect 19794 10792 19800 10804
rect 19755 10764 19800 10792
rect 19794 10752 19800 10764
rect 19852 10752 19858 10804
rect 25590 10792 25596 10804
rect 25240 10764 25596 10792
rect 15488 10724 15516 10752
rect 16482 10724 16488 10736
rect 15488 10696 16488 10724
rect 16482 10684 16488 10696
rect 16540 10684 16546 10736
rect 2866 10616 2872 10668
rect 2924 10656 2930 10668
rect 3970 10656 3976 10668
rect 2924 10628 3976 10656
rect 2924 10616 2930 10628
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 4890 10656 4896 10668
rect 4387 10628 4896 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 8846 10656 8852 10668
rect 8807 10628 8852 10656
rect 8846 10616 8852 10628
rect 8904 10616 8910 10668
rect 9582 10656 9588 10668
rect 9495 10628 9588 10656
rect 9582 10616 9588 10628
rect 9640 10656 9646 10668
rect 10965 10659 11023 10665
rect 10965 10656 10977 10659
rect 9640 10628 10977 10656
rect 9640 10616 9646 10628
rect 10965 10625 10977 10628
rect 11011 10625 11023 10659
rect 13538 10656 13544 10668
rect 10965 10619 11023 10625
rect 13004 10628 13544 10656
rect 3326 10548 3332 10600
rect 3384 10588 3390 10600
rect 3421 10591 3479 10597
rect 3421 10588 3433 10591
rect 3384 10560 3433 10588
rect 3384 10548 3390 10560
rect 3421 10557 3433 10560
rect 3467 10557 3479 10591
rect 3421 10551 3479 10557
rect 8294 10548 8300 10600
rect 8352 10588 8358 10600
rect 9600 10588 9628 10616
rect 8352 10560 9628 10588
rect 9677 10591 9735 10597
rect 8352 10548 8358 10560
rect 9677 10557 9689 10591
rect 9723 10588 9735 10591
rect 9858 10588 9864 10600
rect 9723 10560 9864 10588
rect 9723 10557 9735 10560
rect 9677 10551 9735 10557
rect 9858 10548 9864 10560
rect 9916 10588 9922 10600
rect 10870 10588 10876 10600
rect 9916 10560 10876 10588
rect 9916 10548 9922 10560
rect 10870 10548 10876 10560
rect 10928 10548 10934 10600
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 11514 10588 11520 10600
rect 11112 10560 11520 10588
rect 11112 10548 11118 10560
rect 11514 10548 11520 10560
rect 11572 10548 11578 10600
rect 11882 10548 11888 10600
rect 11940 10588 11946 10600
rect 13004 10597 13032 10628
rect 13538 10616 13544 10628
rect 13596 10656 13602 10668
rect 14918 10656 14924 10668
rect 13596 10628 14924 10656
rect 13596 10616 13602 10628
rect 14918 10616 14924 10628
rect 14976 10616 14982 10668
rect 15473 10659 15531 10665
rect 15473 10625 15485 10659
rect 15519 10656 15531 10659
rect 15654 10656 15660 10668
rect 15519 10628 15660 10656
rect 15519 10625 15531 10628
rect 15473 10619 15531 10625
rect 15654 10616 15660 10628
rect 15712 10616 15718 10668
rect 18414 10656 18420 10668
rect 16408 10628 18420 10656
rect 12253 10591 12311 10597
rect 12253 10588 12265 10591
rect 11940 10560 12265 10588
rect 11940 10548 11946 10560
rect 12253 10557 12265 10560
rect 12299 10557 12311 10591
rect 12253 10551 12311 10557
rect 12989 10591 13047 10597
rect 12989 10557 13001 10591
rect 13035 10557 13047 10591
rect 13262 10588 13268 10600
rect 13223 10560 13268 10588
rect 12989 10551 13047 10557
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 13449 10591 13507 10597
rect 13449 10557 13461 10591
rect 13495 10557 13507 10591
rect 13449 10551 13507 10557
rect 5350 10480 5356 10532
rect 5408 10480 5414 10532
rect 8570 10520 8576 10532
rect 8531 10492 8576 10520
rect 8570 10480 8576 10492
rect 8628 10480 8634 10532
rect 13170 10480 13176 10532
rect 13228 10520 13234 10532
rect 13464 10520 13492 10551
rect 13722 10548 13728 10600
rect 13780 10588 13786 10600
rect 13909 10591 13967 10597
rect 13909 10588 13921 10591
rect 13780 10560 13921 10588
rect 13780 10548 13786 10560
rect 13909 10557 13921 10560
rect 13955 10557 13967 10591
rect 14182 10588 14188 10600
rect 14143 10560 14188 10588
rect 13909 10551 13967 10557
rect 14182 10548 14188 10560
rect 14240 10548 14246 10600
rect 15194 10588 15200 10600
rect 15155 10560 15200 10588
rect 15194 10548 15200 10560
rect 15252 10548 15258 10600
rect 16408 10597 16436 10628
rect 18414 10616 18420 10628
rect 18472 10616 18478 10668
rect 18598 10656 18604 10668
rect 18559 10628 18604 10656
rect 18598 10616 18604 10628
rect 18656 10616 18662 10668
rect 21177 10659 21235 10665
rect 21177 10625 21189 10659
rect 21223 10656 21235 10659
rect 21266 10656 21272 10668
rect 21223 10628 21272 10656
rect 21223 10625 21235 10628
rect 21177 10619 21235 10625
rect 16209 10591 16267 10597
rect 16209 10557 16221 10591
rect 16255 10557 16267 10591
rect 16209 10551 16267 10557
rect 16393 10591 16451 10597
rect 16393 10557 16405 10591
rect 16439 10557 16451 10591
rect 16393 10551 16451 10557
rect 14090 10520 14096 10532
rect 13228 10492 14096 10520
rect 13228 10480 13234 10492
rect 14090 10480 14096 10492
rect 14148 10480 14154 10532
rect 8202 10452 8208 10464
rect 8163 10424 8208 10452
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 8662 10452 8668 10464
rect 8623 10424 8668 10452
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 10226 10412 10232 10464
rect 10284 10452 10290 10464
rect 10781 10455 10839 10461
rect 10781 10452 10793 10455
rect 10284 10424 10793 10452
rect 10284 10412 10290 10424
rect 10781 10421 10793 10424
rect 10827 10421 10839 10455
rect 10781 10415 10839 10421
rect 10873 10455 10931 10461
rect 10873 10421 10885 10455
rect 10919 10452 10931 10455
rect 11054 10452 11060 10464
rect 10919 10424 11060 10452
rect 10919 10421 10931 10424
rect 10873 10415 10931 10421
rect 11054 10412 11060 10424
rect 11112 10412 11118 10464
rect 13262 10412 13268 10464
rect 13320 10452 13326 10464
rect 14001 10455 14059 10461
rect 14001 10452 14013 10455
rect 13320 10424 14013 10452
rect 13320 10412 13326 10424
rect 14001 10421 14013 10424
rect 14047 10421 14059 10455
rect 15470 10452 15476 10464
rect 15431 10424 15476 10452
rect 14001 10415 14059 10421
rect 15470 10412 15476 10424
rect 15528 10412 15534 10464
rect 16224 10452 16252 10551
rect 17218 10548 17224 10600
rect 17276 10588 17282 10600
rect 17589 10591 17647 10597
rect 17589 10588 17601 10591
rect 17276 10560 17601 10588
rect 17276 10548 17282 10560
rect 17589 10557 17601 10560
rect 17635 10557 17647 10591
rect 17589 10551 17647 10557
rect 17865 10591 17923 10597
rect 17865 10557 17877 10591
rect 17911 10557 17923 10591
rect 18230 10588 18236 10600
rect 18191 10560 18236 10588
rect 17865 10551 17923 10557
rect 16301 10523 16359 10529
rect 16301 10489 16313 10523
rect 16347 10520 16359 10523
rect 17880 10520 17908 10551
rect 18230 10548 18236 10560
rect 18288 10548 18294 10600
rect 18693 10591 18751 10597
rect 18693 10557 18705 10591
rect 18739 10557 18751 10591
rect 19242 10588 19248 10600
rect 19203 10560 19248 10588
rect 18693 10551 18751 10557
rect 16347 10492 17908 10520
rect 16347 10489 16359 10492
rect 16301 10483 16359 10489
rect 18138 10480 18144 10532
rect 18196 10520 18202 10532
rect 18708 10520 18736 10551
rect 19242 10548 19248 10560
rect 19300 10548 19306 10600
rect 18196 10492 18736 10520
rect 18196 10480 18202 10492
rect 19978 10480 19984 10532
rect 20036 10520 20042 10532
rect 20910 10523 20968 10529
rect 20910 10520 20922 10523
rect 20036 10492 20922 10520
rect 20036 10480 20042 10492
rect 20910 10489 20922 10492
rect 20956 10489 20968 10523
rect 20910 10483 20968 10489
rect 16390 10452 16396 10464
rect 16224 10424 16396 10452
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 20806 10412 20812 10464
rect 20864 10452 20870 10464
rect 21192 10452 21220 10619
rect 21266 10616 21272 10628
rect 21324 10616 21330 10668
rect 24397 10659 24455 10665
rect 24397 10625 24409 10659
rect 24443 10656 24455 10659
rect 24578 10656 24584 10668
rect 24443 10628 24584 10656
rect 24443 10625 24455 10628
rect 24397 10619 24455 10625
rect 24578 10616 24584 10628
rect 24636 10656 24642 10668
rect 25133 10659 25191 10665
rect 25133 10656 25145 10659
rect 24636 10628 25145 10656
rect 24636 10616 24642 10628
rect 25133 10625 25145 10628
rect 25179 10656 25191 10659
rect 25240 10656 25268 10764
rect 25590 10752 25596 10764
rect 25648 10752 25654 10804
rect 26878 10792 26884 10804
rect 26839 10764 26884 10792
rect 26878 10752 26884 10764
rect 26936 10752 26942 10804
rect 29181 10795 29239 10801
rect 29181 10761 29193 10795
rect 29227 10792 29239 10795
rect 29546 10792 29552 10804
rect 29227 10764 29552 10792
rect 29227 10761 29239 10764
rect 29181 10755 29239 10761
rect 29546 10752 29552 10764
rect 29604 10752 29610 10804
rect 29638 10752 29644 10804
rect 29696 10792 29702 10804
rect 31757 10795 31815 10801
rect 31757 10792 31769 10795
rect 29696 10764 31769 10792
rect 29696 10752 29702 10764
rect 31757 10761 31769 10764
rect 31803 10761 31815 10795
rect 33134 10792 33140 10804
rect 33095 10764 33140 10792
rect 31757 10755 31815 10761
rect 33134 10752 33140 10764
rect 33192 10752 33198 10804
rect 29411 10727 29469 10733
rect 29411 10693 29423 10727
rect 29457 10724 29469 10727
rect 31202 10724 31208 10736
rect 29457 10696 31208 10724
rect 29457 10693 29469 10696
rect 29411 10687 29469 10693
rect 31202 10684 31208 10696
rect 31260 10684 31266 10736
rect 25406 10656 25412 10668
rect 25179 10628 25268 10656
rect 25367 10628 25412 10656
rect 25179 10625 25191 10628
rect 25133 10619 25191 10625
rect 25406 10616 25412 10628
rect 25464 10616 25470 10668
rect 29273 10659 29331 10665
rect 29273 10625 29285 10659
rect 29319 10656 29331 10659
rect 29638 10656 29644 10668
rect 29319 10628 29644 10656
rect 29319 10625 29331 10628
rect 29273 10619 29331 10625
rect 29638 10616 29644 10628
rect 29696 10616 29702 10668
rect 30374 10616 30380 10668
rect 30432 10656 30438 10668
rect 30745 10659 30803 10665
rect 30745 10656 30757 10659
rect 30432 10628 30757 10656
rect 30432 10616 30438 10628
rect 30745 10625 30757 10628
rect 30791 10625 30803 10659
rect 31018 10656 31024 10668
rect 30745 10619 30803 10625
rect 30944 10628 31024 10656
rect 23750 10548 23756 10600
rect 23808 10588 23814 10600
rect 24130 10591 24188 10597
rect 24130 10588 24142 10591
rect 23808 10560 24142 10588
rect 23808 10548 23814 10560
rect 24130 10557 24142 10560
rect 24176 10557 24188 10591
rect 29086 10588 29092 10600
rect 29047 10560 29092 10588
rect 24130 10551 24188 10557
rect 29086 10548 29092 10560
rect 29144 10548 29150 10600
rect 29549 10591 29607 10597
rect 29549 10557 29561 10591
rect 29595 10557 29607 10591
rect 30650 10588 30656 10600
rect 30611 10560 30656 10588
rect 29549 10551 29607 10557
rect 27154 10520 27160 10532
rect 26634 10492 27160 10520
rect 27154 10480 27160 10492
rect 27212 10520 27218 10532
rect 28258 10520 28264 10532
rect 27212 10492 28264 10520
rect 27212 10480 27218 10492
rect 28258 10480 28264 10492
rect 28316 10480 28322 10532
rect 23014 10452 23020 10464
rect 20864 10424 21220 10452
rect 22975 10424 23020 10452
rect 20864 10412 20870 10424
rect 23014 10412 23020 10424
rect 23072 10412 23078 10464
rect 29564 10452 29592 10551
rect 30650 10548 30656 10560
rect 30708 10548 30714 10600
rect 30944 10597 30972 10628
rect 31018 10616 31024 10628
rect 31076 10616 31082 10668
rect 33410 10656 33416 10668
rect 33060 10628 33416 10656
rect 30929 10591 30987 10597
rect 30929 10557 30941 10591
rect 30975 10557 30987 10591
rect 30929 10551 30987 10557
rect 31113 10591 31171 10597
rect 31113 10557 31125 10591
rect 31159 10557 31171 10591
rect 31113 10551 31171 10557
rect 31128 10520 31156 10551
rect 31478 10548 31484 10600
rect 31536 10588 31542 10600
rect 33060 10597 33088 10628
rect 33410 10616 33416 10628
rect 33468 10616 33474 10668
rect 31573 10591 31631 10597
rect 31573 10588 31585 10591
rect 31536 10560 31585 10588
rect 31536 10548 31542 10560
rect 31573 10557 31585 10560
rect 31619 10557 31631 10591
rect 31573 10551 31631 10557
rect 33045 10591 33103 10597
rect 33045 10557 33057 10591
rect 33091 10557 33103 10591
rect 33226 10588 33232 10600
rect 33187 10560 33232 10588
rect 33045 10551 33103 10557
rect 33226 10548 33232 10560
rect 33284 10548 33290 10600
rect 31662 10520 31668 10532
rect 31128 10492 31668 10520
rect 31662 10480 31668 10492
rect 31720 10480 31726 10532
rect 31294 10452 31300 10464
rect 29564 10424 31300 10452
rect 31294 10412 31300 10424
rect 31352 10412 31358 10464
rect 1104 10362 34316 10384
rect 1104 10310 12052 10362
rect 12104 10310 12116 10362
rect 12168 10310 12180 10362
rect 12232 10310 12244 10362
rect 12296 10310 23123 10362
rect 23175 10310 23187 10362
rect 23239 10310 23251 10362
rect 23303 10310 23315 10362
rect 23367 10310 34316 10362
rect 1104 10288 34316 10310
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 10226 10248 10232 10260
rect 2832 10220 2877 10248
rect 10187 10220 10232 10248
rect 2832 10208 2838 10220
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 13262 10248 13268 10260
rect 13223 10220 13268 10248
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 14734 10248 14740 10260
rect 14695 10220 14740 10248
rect 14734 10208 14740 10220
rect 14792 10248 14798 10260
rect 15562 10248 15568 10260
rect 14792 10220 15568 10248
rect 14792 10208 14798 10220
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 16482 10208 16488 10260
rect 16540 10248 16546 10260
rect 19978 10248 19984 10260
rect 16540 10220 19564 10248
rect 19939 10220 19984 10248
rect 16540 10208 16546 10220
rect 7377 10183 7435 10189
rect 7377 10149 7389 10183
rect 7423 10180 7435 10183
rect 8481 10183 8539 10189
rect 8481 10180 8493 10183
rect 7423 10152 8493 10180
rect 7423 10149 7435 10152
rect 7377 10143 7435 10149
rect 8481 10149 8493 10152
rect 8527 10149 8539 10183
rect 9306 10180 9312 10192
rect 8481 10143 8539 10149
rect 8772 10152 9312 10180
rect 8772 10124 8800 10152
rect 9306 10140 9312 10152
rect 9364 10180 9370 10192
rect 9364 10152 10456 10180
rect 9364 10140 9370 10152
rect 8202 10112 8208 10124
rect 8163 10084 8208 10112
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 8297 10115 8355 10121
rect 8297 10081 8309 10115
rect 8343 10112 8355 10115
rect 8754 10112 8760 10124
rect 8343 10084 8760 10112
rect 8343 10081 8355 10084
rect 8297 10075 8355 10081
rect 8754 10072 8760 10084
rect 8812 10072 8818 10124
rect 9398 10072 9404 10124
rect 9456 10112 9462 10124
rect 10428 10121 10456 10152
rect 12802 10140 12808 10192
rect 12860 10180 12866 10192
rect 13633 10183 13691 10189
rect 13633 10180 13645 10183
rect 12860 10152 13645 10180
rect 12860 10140 12866 10152
rect 13633 10149 13645 10152
rect 13679 10149 13691 10183
rect 13633 10143 13691 10149
rect 15470 10140 15476 10192
rect 15528 10180 15534 10192
rect 15850 10183 15908 10189
rect 15850 10180 15862 10183
rect 15528 10152 15862 10180
rect 15528 10140 15534 10152
rect 15850 10149 15862 10152
rect 15896 10149 15908 10183
rect 15850 10143 15908 10149
rect 16758 10140 16764 10192
rect 16816 10180 16822 10192
rect 17310 10180 17316 10192
rect 16816 10152 17316 10180
rect 16816 10140 16822 10152
rect 17310 10140 17316 10152
rect 17368 10180 17374 10192
rect 17368 10152 17816 10180
rect 17368 10140 17374 10152
rect 9493 10115 9551 10121
rect 9493 10112 9505 10115
rect 9456 10084 9505 10112
rect 9456 10072 9462 10084
rect 9493 10081 9505 10084
rect 9539 10081 9551 10115
rect 9493 10075 9551 10081
rect 10413 10115 10471 10121
rect 10413 10081 10425 10115
rect 10459 10081 10471 10115
rect 10413 10075 10471 10081
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10112 10563 10115
rect 11330 10112 11336 10124
rect 10551 10084 11008 10112
rect 11291 10084 11336 10112
rect 10551 10081 10563 10084
rect 10505 10075 10563 10081
rect 2866 10044 2872 10056
rect 2827 10016 2872 10044
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10044 3111 10047
rect 3326 10044 3332 10056
rect 3099 10016 3332 10044
rect 3099 10013 3111 10016
rect 3053 10007 3111 10013
rect 3326 10004 3332 10016
rect 3384 10004 3390 10056
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 7653 10047 7711 10053
rect 7653 10013 7665 10047
rect 7699 10044 7711 10047
rect 8110 10044 8116 10056
rect 7699 10016 8116 10044
rect 7699 10013 7711 10016
rect 7653 10007 7711 10013
rect 7484 9976 7512 10007
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 8481 10047 8539 10053
rect 8481 10013 8493 10047
rect 8527 10044 8539 10047
rect 10134 10044 10140 10056
rect 8527 10016 10140 10044
rect 8527 10013 8539 10016
rect 8481 10007 8539 10013
rect 10134 10004 10140 10016
rect 10192 10044 10198 10056
rect 10229 10047 10287 10053
rect 10229 10044 10241 10047
rect 10192 10016 10241 10044
rect 10192 10004 10198 10016
rect 10229 10013 10241 10016
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 8386 9976 8392 9988
rect 7484 9948 8392 9976
rect 8386 9936 8392 9948
rect 8444 9936 8450 9988
rect 10980 9985 11008 10084
rect 11330 10072 11336 10084
rect 11388 10072 11394 10124
rect 12897 10115 12955 10121
rect 12897 10081 12909 10115
rect 12943 10081 12955 10115
rect 13446 10112 13452 10124
rect 13407 10084 13452 10112
rect 12897 10075 12955 10081
rect 11422 10044 11428 10056
rect 11383 10016 11428 10044
rect 11422 10004 11428 10016
rect 11480 10004 11486 10056
rect 11514 10004 11520 10056
rect 11572 10044 11578 10056
rect 11572 10016 11617 10044
rect 11572 10004 11578 10016
rect 10965 9979 11023 9985
rect 10965 9945 10977 9979
rect 11011 9945 11023 9979
rect 10965 9939 11023 9945
rect 1762 9868 1768 9920
rect 1820 9908 1826 9920
rect 2409 9911 2467 9917
rect 2409 9908 2421 9911
rect 1820 9880 2421 9908
rect 1820 9868 1826 9880
rect 2409 9877 2421 9880
rect 2455 9877 2467 9911
rect 2409 9871 2467 9877
rect 7009 9911 7067 9917
rect 7009 9877 7021 9911
rect 7055 9908 7067 9911
rect 7098 9908 7104 9920
rect 7055 9880 7104 9908
rect 7055 9877 7067 9880
rect 7009 9871 7067 9877
rect 7098 9868 7104 9880
rect 7156 9868 7162 9920
rect 9585 9911 9643 9917
rect 9585 9877 9597 9911
rect 9631 9908 9643 9911
rect 9674 9908 9680 9920
rect 9631 9880 9680 9908
rect 9631 9877 9643 9880
rect 9585 9871 9643 9877
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 11882 9868 11888 9920
rect 11940 9908 11946 9920
rect 12713 9911 12771 9917
rect 12713 9908 12725 9911
rect 11940 9880 12725 9908
rect 11940 9868 11946 9880
rect 12713 9877 12725 9880
rect 12759 9877 12771 9911
rect 12912 9908 12940 10075
rect 13446 10072 13452 10084
rect 13504 10072 13510 10124
rect 16114 10112 16120 10124
rect 16075 10084 16120 10112
rect 16114 10072 16120 10084
rect 16172 10072 16178 10124
rect 16666 10112 16672 10124
rect 16627 10084 16672 10112
rect 16666 10072 16672 10084
rect 16724 10072 16730 10124
rect 16942 10112 16948 10124
rect 16903 10084 16948 10112
rect 16942 10072 16948 10084
rect 17000 10072 17006 10124
rect 17402 10112 17408 10124
rect 17363 10084 17408 10112
rect 17402 10072 17408 10084
rect 17460 10072 17466 10124
rect 17788 10121 17816 10152
rect 17773 10115 17831 10121
rect 17773 10081 17785 10115
rect 17819 10081 17831 10115
rect 17773 10075 17831 10081
rect 17954 10072 17960 10124
rect 18012 10112 18018 10124
rect 18141 10115 18199 10121
rect 18141 10112 18153 10115
rect 18012 10084 18153 10112
rect 18012 10072 18018 10084
rect 18141 10081 18153 10084
rect 18187 10081 18199 10115
rect 19536 10112 19564 10220
rect 19978 10208 19984 10220
rect 20036 10208 20042 10260
rect 22189 10251 22247 10257
rect 22189 10217 22201 10251
rect 22235 10248 22247 10251
rect 22554 10248 22560 10260
rect 22235 10220 22560 10248
rect 22235 10217 22247 10220
rect 22189 10211 22247 10217
rect 22554 10208 22560 10220
rect 22612 10208 22618 10260
rect 23842 10208 23848 10260
rect 23900 10248 23906 10260
rect 23937 10251 23995 10257
rect 23937 10248 23949 10251
rect 23900 10220 23949 10248
rect 23900 10208 23906 10220
rect 23937 10217 23949 10220
rect 23983 10217 23995 10251
rect 23937 10211 23995 10217
rect 29638 10208 29644 10260
rect 29696 10248 29702 10260
rect 29696 10220 31708 10248
rect 29696 10208 29702 10220
rect 23201 10183 23259 10189
rect 23201 10180 23213 10183
rect 20272 10152 23213 10180
rect 20272 10121 20300 10152
rect 23201 10149 23213 10152
rect 23247 10149 23259 10183
rect 23201 10143 23259 10149
rect 27154 10140 27160 10192
rect 27212 10180 27218 10192
rect 27212 10152 27370 10180
rect 27212 10140 27218 10152
rect 30190 10140 30196 10192
rect 30248 10180 30254 10192
rect 30248 10152 30972 10180
rect 30248 10140 30254 10152
rect 20165 10115 20223 10121
rect 20165 10112 20177 10115
rect 19536 10084 20177 10112
rect 18141 10075 18199 10081
rect 20165 10081 20177 10084
rect 20211 10081 20223 10115
rect 20165 10075 20223 10081
rect 20257 10115 20315 10121
rect 20257 10081 20269 10115
rect 20303 10081 20315 10115
rect 20806 10112 20812 10124
rect 20767 10084 20812 10112
rect 20257 10075 20315 10081
rect 17310 10004 17316 10056
rect 17368 10044 17374 10056
rect 17681 10047 17739 10053
rect 17681 10044 17693 10047
rect 17368 10016 17693 10044
rect 17368 10004 17374 10016
rect 17681 10013 17693 10016
rect 17727 10013 17739 10047
rect 19978 10044 19984 10056
rect 19939 10016 19984 10044
rect 17681 10007 17739 10013
rect 19978 10004 19984 10016
rect 20036 10004 20042 10056
rect 20180 10044 20208 10075
rect 20806 10072 20812 10084
rect 20864 10072 20870 10124
rect 21076 10115 21134 10121
rect 21076 10081 21088 10115
rect 21122 10112 21134 10115
rect 21358 10112 21364 10124
rect 21122 10084 21364 10112
rect 21122 10081 21134 10084
rect 21076 10075 21134 10081
rect 21358 10072 21364 10084
rect 21416 10072 21422 10124
rect 22649 10115 22707 10121
rect 22649 10112 22661 10115
rect 22066 10084 22661 10112
rect 20530 10044 20536 10056
rect 20180 10016 20536 10044
rect 20530 10004 20536 10016
rect 20588 10004 20594 10056
rect 17144 9948 20300 9976
rect 17144 9920 17172 9948
rect 17126 9908 17132 9920
rect 12912 9880 17132 9908
rect 12713 9871 12771 9877
rect 17126 9868 17132 9880
rect 17184 9868 17190 9920
rect 20272 9908 20300 9948
rect 22066 9908 22094 10084
rect 22649 10081 22661 10084
rect 22695 10081 22707 10115
rect 22649 10075 22707 10081
rect 23014 10072 23020 10124
rect 23072 10112 23078 10124
rect 23293 10115 23351 10121
rect 23293 10112 23305 10115
rect 23072 10084 23305 10112
rect 23072 10072 23078 10084
rect 23293 10081 23305 10084
rect 23339 10112 23351 10115
rect 23845 10115 23903 10121
rect 23845 10112 23857 10115
rect 23339 10084 23857 10112
rect 23339 10081 23351 10084
rect 23293 10075 23351 10081
rect 23845 10081 23857 10084
rect 23891 10081 23903 10115
rect 23845 10075 23903 10081
rect 24029 10115 24087 10121
rect 24029 10081 24041 10115
rect 24075 10081 24087 10115
rect 24029 10075 24087 10081
rect 22370 10004 22376 10056
rect 22428 10044 22434 10056
rect 24044 10044 24072 10075
rect 25590 10072 25596 10124
rect 25648 10112 25654 10124
rect 26605 10115 26663 10121
rect 26605 10112 26617 10115
rect 25648 10084 26617 10112
rect 25648 10072 25654 10084
rect 26605 10081 26617 10084
rect 26651 10081 26663 10115
rect 30742 10112 30748 10124
rect 30703 10084 30748 10112
rect 26605 10075 26663 10081
rect 30742 10072 30748 10084
rect 30800 10072 30806 10124
rect 30944 10121 30972 10152
rect 30837 10115 30895 10121
rect 30837 10081 30849 10115
rect 30883 10081 30895 10115
rect 30837 10075 30895 10081
rect 30929 10115 30987 10121
rect 30929 10081 30941 10115
rect 30975 10081 30987 10115
rect 31110 10112 31116 10124
rect 31071 10084 31116 10112
rect 30929 10075 30987 10081
rect 22428 10016 24072 10044
rect 26881 10047 26939 10053
rect 22428 10004 22434 10016
rect 26881 10013 26893 10047
rect 26927 10044 26939 10047
rect 30469 10047 30527 10053
rect 30469 10044 30481 10047
rect 26927 10016 30481 10044
rect 26927 10013 26939 10016
rect 26881 10007 26939 10013
rect 30469 10013 30481 10016
rect 30515 10013 30527 10047
rect 30469 10007 30527 10013
rect 29086 9936 29092 9988
rect 29144 9976 29150 9988
rect 30852 9976 30880 10075
rect 31110 10072 31116 10084
rect 31168 10112 31174 10124
rect 31478 10112 31484 10124
rect 31168 10084 31484 10112
rect 31168 10072 31174 10084
rect 31478 10072 31484 10084
rect 31536 10072 31542 10124
rect 31573 10115 31631 10121
rect 31573 10081 31585 10115
rect 31619 10081 31631 10115
rect 31680 10112 31708 10220
rect 32306 10140 32312 10192
rect 32364 10180 32370 10192
rect 32585 10183 32643 10189
rect 32585 10180 32597 10183
rect 32364 10152 32597 10180
rect 32364 10140 32370 10152
rect 32585 10149 32597 10152
rect 32631 10180 32643 10183
rect 32631 10152 33456 10180
rect 32631 10149 32643 10152
rect 32585 10143 32643 10149
rect 31757 10115 31815 10121
rect 31757 10112 31769 10115
rect 31680 10084 31769 10112
rect 31573 10075 31631 10081
rect 31757 10081 31769 10084
rect 31803 10081 31815 10115
rect 32398 10112 32404 10124
rect 32359 10084 32404 10112
rect 31757 10075 31815 10081
rect 31294 10004 31300 10056
rect 31352 10044 31358 10056
rect 31588 10044 31616 10075
rect 31352 10016 31616 10044
rect 31772 10044 31800 10075
rect 32398 10072 32404 10084
rect 32456 10072 32462 10124
rect 33428 10121 33456 10152
rect 33229 10115 33287 10121
rect 33229 10081 33241 10115
rect 33275 10081 33287 10115
rect 33229 10075 33287 10081
rect 33413 10115 33471 10121
rect 33413 10081 33425 10115
rect 33459 10081 33471 10115
rect 33413 10075 33471 10081
rect 33244 10044 33272 10075
rect 31772 10016 33272 10044
rect 31352 10004 31358 10016
rect 29144 9948 30880 9976
rect 29144 9936 29150 9948
rect 31662 9936 31668 9988
rect 31720 9976 31726 9988
rect 31849 9979 31907 9985
rect 31849 9976 31861 9979
rect 31720 9948 31861 9976
rect 31720 9936 31726 9948
rect 31849 9945 31861 9948
rect 31895 9945 31907 9979
rect 33244 9976 33272 10016
rect 33410 9976 33416 9988
rect 33244 9948 33416 9976
rect 31849 9939 31907 9945
rect 33410 9936 33416 9948
rect 33468 9936 33474 9988
rect 22830 9908 22836 9920
rect 20272 9880 22094 9908
rect 22791 9880 22836 9908
rect 22830 9868 22836 9880
rect 22888 9868 22894 9920
rect 28350 9908 28356 9920
rect 28311 9880 28356 9908
rect 28350 9868 28356 9880
rect 28408 9868 28414 9920
rect 32769 9911 32827 9917
rect 32769 9877 32781 9911
rect 32815 9908 32827 9911
rect 33134 9908 33140 9920
rect 32815 9880 33140 9908
rect 32815 9877 32827 9880
rect 32769 9871 32827 9877
rect 33134 9868 33140 9880
rect 33192 9868 33198 9920
rect 33318 9908 33324 9920
rect 33279 9880 33324 9908
rect 33318 9868 33324 9880
rect 33376 9868 33382 9920
rect 1104 9818 34316 9840
rect 1104 9766 6517 9818
rect 6569 9766 6581 9818
rect 6633 9766 6645 9818
rect 6697 9766 6709 9818
rect 6761 9766 17588 9818
rect 17640 9766 17652 9818
rect 17704 9766 17716 9818
rect 17768 9766 17780 9818
rect 17832 9766 28658 9818
rect 28710 9766 28722 9818
rect 28774 9766 28786 9818
rect 28838 9766 28850 9818
rect 28902 9766 34316 9818
rect 1104 9744 34316 9766
rect 2866 9664 2872 9716
rect 2924 9704 2930 9716
rect 3191 9707 3249 9713
rect 3191 9704 3203 9707
rect 2924 9676 3203 9704
rect 2924 9664 2930 9676
rect 3191 9673 3203 9676
rect 3237 9673 3249 9707
rect 3191 9667 3249 9673
rect 8570 9664 8576 9716
rect 8628 9704 8634 9716
rect 9125 9707 9183 9713
rect 9125 9704 9137 9707
rect 8628 9676 9137 9704
rect 8628 9664 8634 9676
rect 9125 9673 9137 9676
rect 9171 9673 9183 9707
rect 9125 9667 9183 9673
rect 11330 9664 11336 9716
rect 11388 9704 11394 9716
rect 12069 9707 12127 9713
rect 12069 9704 12081 9707
rect 11388 9676 12081 9704
rect 11388 9664 11394 9676
rect 12069 9673 12081 9676
rect 12115 9673 12127 9707
rect 15654 9704 15660 9716
rect 15615 9676 15660 9704
rect 12069 9667 12127 9673
rect 15654 9664 15660 9676
rect 15712 9664 15718 9716
rect 19797 9707 19855 9713
rect 19797 9673 19809 9707
rect 19843 9704 19855 9707
rect 19978 9704 19984 9716
rect 19843 9676 19984 9704
rect 19843 9673 19855 9676
rect 19797 9667 19855 9673
rect 19978 9664 19984 9676
rect 20036 9664 20042 9716
rect 21358 9704 21364 9716
rect 21319 9676 21364 9704
rect 21358 9664 21364 9676
rect 21416 9664 21422 9716
rect 29917 9707 29975 9713
rect 29917 9673 29929 9707
rect 29963 9704 29975 9707
rect 33229 9707 33287 9713
rect 29963 9676 30420 9704
rect 29963 9673 29975 9676
rect 29917 9667 29975 9673
rect 11054 9636 11060 9648
rect 11015 9608 11060 9636
rect 11054 9596 11060 9608
rect 11112 9596 11118 9648
rect 16850 9596 16856 9648
rect 16908 9636 16914 9648
rect 17589 9639 17647 9645
rect 17589 9636 17601 9639
rect 16908 9608 17601 9636
rect 16908 9596 16914 9608
rect 17589 9605 17601 9608
rect 17635 9605 17647 9639
rect 17589 9599 17647 9605
rect 21174 9596 21180 9648
rect 21232 9636 21238 9648
rect 21453 9639 21511 9645
rect 21453 9636 21465 9639
rect 21232 9608 21465 9636
rect 21232 9596 21238 9608
rect 21453 9605 21465 9608
rect 21499 9605 21511 9639
rect 25958 9636 25964 9648
rect 25919 9608 25964 9636
rect 21453 9599 21511 9605
rect 25958 9596 25964 9608
rect 26016 9596 26022 9648
rect 1762 9568 1768 9580
rect 1723 9540 1768 9568
rect 1762 9528 1768 9540
rect 1820 9528 1826 9580
rect 5258 9528 5264 9580
rect 5316 9568 5322 9580
rect 5537 9571 5595 9577
rect 5537 9568 5549 9571
rect 5316 9540 5549 9568
rect 5316 9528 5322 9540
rect 5537 9537 5549 9540
rect 5583 9537 5595 9571
rect 5537 9531 5595 9537
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9537 5687 9571
rect 7098 9568 7104 9580
rect 7059 9540 7104 9568
rect 5629 9531 5687 9537
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1486 9500 1492 9512
rect 1443 9472 1492 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1486 9460 1492 9472
rect 1544 9460 1550 9512
rect 3786 9460 3792 9512
rect 3844 9500 3850 9512
rect 3881 9503 3939 9509
rect 3881 9500 3893 9503
rect 3844 9472 3893 9500
rect 3844 9460 3850 9472
rect 3881 9469 3893 9472
rect 3927 9469 3939 9503
rect 3881 9463 3939 9469
rect 4430 9460 4436 9512
rect 4488 9500 4494 9512
rect 5644 9500 5672 9531
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 8573 9571 8631 9577
rect 8573 9537 8585 9571
rect 8619 9568 8631 9571
rect 9214 9568 9220 9580
rect 8619 9540 9220 9568
rect 8619 9537 8631 9540
rect 8573 9531 8631 9537
rect 9214 9528 9220 9540
rect 9272 9568 9278 9580
rect 9398 9568 9404 9580
rect 9272 9540 9404 9568
rect 9272 9528 9278 9540
rect 9398 9528 9404 9540
rect 9456 9528 9462 9580
rect 9766 9568 9772 9580
rect 9727 9540 9772 9568
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 12713 9571 12771 9577
rect 12713 9537 12725 9571
rect 12759 9568 12771 9571
rect 12894 9568 12900 9580
rect 12759 9540 12900 9568
rect 12759 9537 12771 9540
rect 12713 9531 12771 9537
rect 12894 9528 12900 9540
rect 12952 9528 12958 9580
rect 13354 9528 13360 9580
rect 13412 9568 13418 9580
rect 13630 9568 13636 9580
rect 13412 9540 13636 9568
rect 13412 9528 13418 9540
rect 13630 9528 13636 9540
rect 13688 9568 13694 9580
rect 13817 9571 13875 9577
rect 13817 9568 13829 9571
rect 13688 9540 13829 9568
rect 13688 9528 13694 9540
rect 13817 9537 13829 9540
rect 13863 9537 13875 9571
rect 13817 9531 13875 9537
rect 21269 9571 21327 9577
rect 21269 9537 21281 9571
rect 21315 9568 21327 9571
rect 21910 9568 21916 9580
rect 21315 9540 21916 9568
rect 21315 9537 21327 9540
rect 21269 9531 21327 9537
rect 21910 9528 21916 9540
rect 21968 9528 21974 9580
rect 24578 9568 24584 9580
rect 24539 9540 24584 9568
rect 24578 9528 24584 9540
rect 24636 9528 24642 9580
rect 6822 9500 6828 9512
rect 4488 9472 5672 9500
rect 6783 9472 6828 9500
rect 4488 9460 4494 9472
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 8662 9460 8668 9512
rect 8720 9500 8726 9512
rect 9490 9500 9496 9512
rect 8720 9472 9496 9500
rect 8720 9460 8726 9472
rect 9490 9460 9496 9472
rect 9548 9500 9554 9512
rect 10321 9503 10379 9509
rect 10321 9500 10333 9503
rect 9548 9472 10333 9500
rect 9548 9460 9554 9472
rect 10321 9469 10333 9472
rect 10367 9469 10379 9503
rect 10321 9463 10379 9469
rect 11149 9503 11207 9509
rect 11149 9469 11161 9503
rect 11195 9469 11207 9503
rect 11149 9463 11207 9469
rect 2314 9392 2320 9444
rect 2372 9392 2378 9444
rect 3326 9392 3332 9444
rect 3384 9432 3390 9444
rect 3697 9435 3755 9441
rect 3697 9432 3709 9435
rect 3384 9404 3709 9432
rect 3384 9392 3390 9404
rect 3697 9401 3709 9404
rect 3743 9401 3755 9435
rect 3697 9395 3755 9401
rect 5445 9435 5503 9441
rect 5445 9401 5457 9435
rect 5491 9432 5503 9435
rect 5626 9432 5632 9444
rect 5491 9404 5632 9432
rect 5491 9401 5503 9404
rect 5445 9395 5503 9401
rect 5626 9392 5632 9404
rect 5684 9392 5690 9444
rect 8110 9392 8116 9444
rect 8168 9392 8174 9444
rect 8386 9392 8392 9444
rect 8444 9432 8450 9444
rect 10413 9435 10471 9441
rect 10413 9432 10425 9435
rect 8444 9404 10425 9432
rect 8444 9392 8450 9404
rect 10413 9401 10425 9404
rect 10459 9401 10471 9435
rect 11164 9432 11192 9463
rect 13446 9460 13452 9512
rect 13504 9500 13510 9512
rect 14461 9503 14519 9509
rect 14461 9500 14473 9503
rect 13504 9472 14473 9500
rect 13504 9460 13510 9472
rect 14461 9469 14473 9472
rect 14507 9469 14519 9503
rect 15562 9500 15568 9512
rect 15523 9472 15568 9500
rect 14461 9463 14519 9469
rect 15562 9460 15568 9472
rect 15620 9460 15626 9512
rect 15749 9503 15807 9509
rect 15749 9469 15761 9503
rect 15795 9500 15807 9503
rect 15838 9500 15844 9512
rect 15795 9472 15844 9500
rect 15795 9469 15807 9472
rect 15749 9463 15807 9469
rect 11422 9432 11428 9444
rect 11164 9404 11428 9432
rect 10413 9395 10471 9401
rect 11422 9392 11428 9404
rect 11480 9432 11486 9444
rect 12437 9435 12495 9441
rect 12437 9432 12449 9435
rect 11480 9404 12449 9432
rect 11480 9392 11486 9404
rect 12437 9401 12449 9404
rect 12483 9432 12495 9435
rect 15764 9432 15792 9463
rect 15838 9460 15844 9472
rect 15896 9460 15902 9512
rect 17310 9500 17316 9512
rect 17271 9472 17316 9500
rect 17310 9460 17316 9472
rect 17368 9460 17374 9512
rect 17589 9503 17647 9509
rect 17589 9469 17601 9503
rect 17635 9500 17647 9503
rect 18598 9500 18604 9512
rect 17635 9472 18604 9500
rect 17635 9469 17647 9472
rect 17589 9463 17647 9469
rect 18598 9460 18604 9472
rect 18656 9460 18662 9512
rect 19705 9503 19763 9509
rect 19705 9469 19717 9503
rect 19751 9500 19763 9503
rect 19794 9500 19800 9512
rect 19751 9472 19800 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 19794 9460 19800 9472
rect 19852 9460 19858 9512
rect 19889 9503 19947 9509
rect 19889 9469 19901 9503
rect 19935 9469 19947 9503
rect 19889 9463 19947 9469
rect 19904 9432 19932 9463
rect 20346 9460 20352 9512
rect 20404 9500 20410 9512
rect 20625 9503 20683 9509
rect 20625 9500 20637 9503
rect 20404 9472 20637 9500
rect 20404 9460 20410 9472
rect 20625 9469 20637 9472
rect 20671 9469 20683 9503
rect 21542 9500 21548 9512
rect 21503 9472 21548 9500
rect 20625 9463 20683 9469
rect 21542 9460 21548 9472
rect 21600 9460 21606 9512
rect 22554 9500 22560 9512
rect 22515 9472 22560 9500
rect 22554 9460 22560 9472
rect 22612 9460 22618 9512
rect 23845 9503 23903 9509
rect 23845 9469 23857 9503
rect 23891 9500 23903 9503
rect 24394 9500 24400 9512
rect 23891 9472 24400 9500
rect 23891 9469 23903 9472
rect 23845 9463 23903 9469
rect 24394 9460 24400 9472
rect 24452 9460 24458 9512
rect 28994 9500 29000 9512
rect 28955 9472 29000 9500
rect 28994 9460 29000 9472
rect 29052 9460 29058 9512
rect 29454 9500 29460 9512
rect 29415 9472 29460 9500
rect 29454 9460 29460 9472
rect 29512 9460 29518 9512
rect 29730 9500 29736 9512
rect 29691 9472 29736 9500
rect 29730 9460 29736 9472
rect 29788 9460 29794 9512
rect 20070 9432 20076 9444
rect 12483 9404 13308 9432
rect 15764 9404 20076 9432
rect 12483 9401 12495 9404
rect 12437 9395 12495 9401
rect 4614 9324 4620 9376
rect 4672 9364 4678 9376
rect 5077 9367 5135 9373
rect 5077 9364 5089 9367
rect 4672 9336 5089 9364
rect 4672 9324 4678 9336
rect 5077 9333 5089 9336
rect 5123 9333 5135 9367
rect 5077 9327 5135 9333
rect 9582 9324 9588 9376
rect 9640 9364 9646 9376
rect 12526 9364 12532 9376
rect 9640 9336 9685 9364
rect 12487 9336 12532 9364
rect 9640 9324 9646 9336
rect 12526 9324 12532 9336
rect 12584 9324 12590 9376
rect 13280 9373 13308 9404
rect 20070 9392 20076 9404
rect 20128 9432 20134 9444
rect 20128 9404 20668 9432
rect 20128 9392 20134 9404
rect 20640 9376 20668 9404
rect 23566 9392 23572 9444
rect 23624 9432 23630 9444
rect 24826 9435 24884 9441
rect 24826 9432 24838 9435
rect 23624 9404 24838 9432
rect 23624 9392 23630 9404
rect 24826 9401 24838 9404
rect 24872 9401 24884 9435
rect 30392 9432 30420 9676
rect 33229 9673 33241 9707
rect 33275 9704 33287 9707
rect 33410 9704 33416 9716
rect 33275 9676 33416 9704
rect 33275 9673 33287 9676
rect 33229 9667 33287 9673
rect 33410 9664 33416 9676
rect 33468 9664 33474 9716
rect 30742 9596 30748 9648
rect 30800 9636 30806 9648
rect 30800 9608 30845 9636
rect 30800 9596 30806 9608
rect 32398 9568 32404 9580
rect 30852 9540 32404 9568
rect 30742 9460 30748 9512
rect 30800 9500 30806 9512
rect 30852 9509 30880 9540
rect 32398 9528 32404 9540
rect 32456 9528 32462 9580
rect 30837 9503 30895 9509
rect 30837 9500 30849 9503
rect 30800 9472 30849 9500
rect 30800 9460 30806 9472
rect 30837 9469 30849 9472
rect 30883 9469 30895 9503
rect 31202 9500 31208 9512
rect 31163 9472 31208 9500
rect 30837 9463 30895 9469
rect 31202 9460 31208 9472
rect 31260 9460 31266 9512
rect 31294 9460 31300 9512
rect 31352 9500 31358 9512
rect 31389 9503 31447 9509
rect 31389 9500 31401 9503
rect 31352 9472 31401 9500
rect 31352 9460 31358 9472
rect 31389 9469 31401 9472
rect 31435 9469 31447 9503
rect 32416 9500 32444 9528
rect 33045 9503 33103 9509
rect 33045 9500 33057 9503
rect 32416 9472 33057 9500
rect 31389 9463 31447 9469
rect 33045 9469 33057 9472
rect 33091 9469 33103 9503
rect 33045 9463 33103 9469
rect 31220 9432 31248 9460
rect 30392 9404 31248 9432
rect 24826 9395 24884 9401
rect 13265 9367 13323 9373
rect 13265 9333 13277 9367
rect 13311 9333 13323 9367
rect 13630 9364 13636 9376
rect 13591 9336 13636 9364
rect 13265 9327 13323 9333
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 13725 9367 13783 9373
rect 13725 9333 13737 9367
rect 13771 9364 13783 9367
rect 14553 9367 14611 9373
rect 14553 9364 14565 9367
rect 13771 9336 14565 9364
rect 13771 9333 13783 9336
rect 13725 9327 13783 9333
rect 14553 9333 14565 9336
rect 14599 9333 14611 9367
rect 14553 9327 14611 9333
rect 20622 9324 20628 9376
rect 20680 9324 20686 9376
rect 20806 9364 20812 9376
rect 20767 9336 20812 9364
rect 20806 9324 20812 9336
rect 20864 9324 20870 9376
rect 20898 9324 20904 9376
rect 20956 9364 20962 9376
rect 22649 9367 22707 9373
rect 22649 9364 22661 9367
rect 20956 9336 22661 9364
rect 20956 9324 20962 9336
rect 22649 9333 22661 9336
rect 22695 9333 22707 9367
rect 22649 9327 22707 9333
rect 23753 9367 23811 9373
rect 23753 9333 23765 9367
rect 23799 9364 23811 9367
rect 23842 9364 23848 9376
rect 23799 9336 23848 9364
rect 23799 9333 23811 9336
rect 23753 9327 23811 9333
rect 23842 9324 23848 9336
rect 23900 9324 23906 9376
rect 1104 9274 34316 9296
rect 1104 9222 12052 9274
rect 12104 9222 12116 9274
rect 12168 9222 12180 9274
rect 12232 9222 12244 9274
rect 12296 9222 23123 9274
rect 23175 9222 23187 9274
rect 23239 9222 23251 9274
rect 23303 9222 23315 9274
rect 23367 9222 34316 9274
rect 1104 9200 34316 9222
rect 5258 9120 5264 9172
rect 5316 9160 5322 9172
rect 6043 9163 6101 9169
rect 6043 9160 6055 9163
rect 5316 9132 6055 9160
rect 5316 9120 5322 9132
rect 6043 9129 6055 9132
rect 6089 9129 6101 9163
rect 6043 9123 6101 9129
rect 8481 9163 8539 9169
rect 8481 9129 8493 9163
rect 8527 9160 8539 9163
rect 9582 9160 9588 9172
rect 8527 9132 9588 9160
rect 8527 9129 8539 9132
rect 8481 9123 8539 9129
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 11425 9163 11483 9169
rect 11425 9129 11437 9163
rect 11471 9160 11483 9163
rect 12526 9160 12532 9172
rect 11471 9132 12532 9160
rect 11471 9129 11483 9132
rect 11425 9123 11483 9129
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 13446 9160 13452 9172
rect 12636 9132 13452 9160
rect 5350 9052 5356 9104
rect 5408 9052 5414 9104
rect 9858 9092 9864 9104
rect 9508 9064 9864 9092
rect 2777 9027 2835 9033
rect 2777 8993 2789 9027
rect 2823 9024 2835 9027
rect 2866 9024 2872 9036
rect 2823 8996 2872 9024
rect 2823 8993 2835 8996
rect 2777 8987 2835 8993
rect 2866 8984 2872 8996
rect 2924 8984 2930 9036
rect 4614 9024 4620 9036
rect 4575 8996 4620 9024
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 8386 9024 8392 9036
rect 8347 8996 8392 9024
rect 8386 8984 8392 8996
rect 8444 8984 8450 9036
rect 9508 9033 9536 9064
rect 9858 9052 9864 9064
rect 9916 9052 9922 9104
rect 10704 9064 11560 9092
rect 8573 9027 8631 9033
rect 8573 8993 8585 9027
rect 8619 8993 8631 9027
rect 8573 8987 8631 8993
rect 9493 9027 9551 9033
rect 9493 8993 9505 9027
rect 9539 8993 9551 9027
rect 9674 9024 9680 9036
rect 9635 8996 9680 9024
rect 9493 8987 9551 8993
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8956 2743 8959
rect 2958 8956 2964 8968
rect 2731 8928 2964 8956
rect 2731 8925 2743 8928
rect 2685 8919 2743 8925
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 4522 8956 4528 8968
rect 4295 8928 4528 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 4522 8916 4528 8928
rect 4580 8916 4586 8968
rect 8588 8956 8616 8987
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 10226 8984 10232 9036
rect 10284 9024 10290 9036
rect 10704 9033 10732 9064
rect 10505 9027 10563 9033
rect 10505 9024 10517 9027
rect 10284 8996 10517 9024
rect 10284 8984 10290 8996
rect 10505 8993 10517 8996
rect 10551 8993 10563 9027
rect 10505 8987 10563 8993
rect 10689 9027 10747 9033
rect 10689 8993 10701 9027
rect 10735 8993 10747 9027
rect 10689 8987 10747 8993
rect 9030 8956 9036 8968
rect 8588 8928 9036 8956
rect 9030 8916 9036 8928
rect 9088 8956 9094 8968
rect 10704 8956 10732 8987
rect 11054 8984 11060 9036
rect 11112 9024 11118 9036
rect 11532 9033 11560 9064
rect 11333 9027 11391 9033
rect 11333 9024 11345 9027
rect 11112 8996 11345 9024
rect 11112 8984 11118 8996
rect 11333 8993 11345 8996
rect 11379 8993 11391 9027
rect 11333 8987 11391 8993
rect 11517 9027 11575 9033
rect 11517 8993 11529 9027
rect 11563 9024 11575 9027
rect 11606 9024 11612 9036
rect 11563 8996 11612 9024
rect 11563 8993 11575 8996
rect 11517 8987 11575 8993
rect 11606 8984 11612 8996
rect 11664 8984 11670 9036
rect 12636 9033 12664 9132
rect 13446 9120 13452 9132
rect 13504 9120 13510 9172
rect 13630 9160 13636 9172
rect 13591 9132 13636 9160
rect 13630 9120 13636 9132
rect 13688 9120 13694 9172
rect 15194 9120 15200 9172
rect 15252 9160 15258 9172
rect 15749 9163 15807 9169
rect 15749 9160 15761 9163
rect 15252 9132 15761 9160
rect 15252 9120 15258 9132
rect 15749 9129 15761 9132
rect 15795 9129 15807 9163
rect 15749 9123 15807 9129
rect 16485 9163 16543 9169
rect 16485 9129 16497 9163
rect 16531 9160 16543 9163
rect 16666 9160 16672 9172
rect 16531 9132 16672 9160
rect 16531 9129 16543 9132
rect 16485 9123 16543 9129
rect 12713 9095 12771 9101
rect 12713 9061 12725 9095
rect 12759 9092 12771 9095
rect 15764 9092 15792 9123
rect 16666 9120 16672 9132
rect 16724 9120 16730 9172
rect 17218 9160 17224 9172
rect 17179 9132 17224 9160
rect 17218 9120 17224 9132
rect 17276 9120 17282 9172
rect 18230 9160 18236 9172
rect 18191 9132 18236 9160
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 20346 9120 20352 9172
rect 20404 9160 20410 9172
rect 21545 9163 21603 9169
rect 20404 9132 21496 9160
rect 20404 9120 20410 9132
rect 20898 9092 20904 9104
rect 12759 9064 13492 9092
rect 15764 9064 16528 9092
rect 12759 9061 12771 9064
rect 12713 9055 12771 9061
rect 12621 9027 12679 9033
rect 12621 8993 12633 9027
rect 12667 8993 12679 9027
rect 12802 9024 12808 9036
rect 12763 8996 12808 9024
rect 12621 8987 12679 8993
rect 12802 8984 12808 8996
rect 12860 8984 12866 9036
rect 13262 9024 13268 9036
rect 13223 8996 13268 9024
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 13464 9033 13492 9064
rect 13449 9027 13507 9033
rect 13449 8993 13461 9027
rect 13495 8993 13507 9027
rect 13449 8987 13507 8993
rect 15841 9027 15899 9033
rect 15841 8993 15853 9027
rect 15887 9024 15899 9027
rect 16114 9024 16120 9036
rect 15887 8996 16120 9024
rect 15887 8993 15899 8996
rect 15841 8987 15899 8993
rect 16114 8984 16120 8996
rect 16172 8984 16178 9036
rect 16206 8984 16212 9036
rect 16264 9024 16270 9036
rect 16500 9033 16528 9064
rect 18800 9064 20904 9092
rect 16301 9027 16359 9033
rect 16301 9024 16313 9027
rect 16264 8996 16313 9024
rect 16264 8984 16270 8996
rect 16301 8993 16313 8996
rect 16347 8993 16359 9027
rect 16301 8987 16359 8993
rect 16485 9027 16543 9033
rect 16485 8993 16497 9027
rect 16531 8993 16543 9027
rect 16485 8987 16543 8993
rect 17129 9027 17187 9033
rect 17129 8993 17141 9027
rect 17175 8993 17187 9027
rect 17129 8987 17187 8993
rect 9088 8928 10732 8956
rect 17144 8956 17172 8987
rect 17218 8984 17224 9036
rect 17276 9024 17282 9036
rect 17313 9027 17371 9033
rect 17313 9024 17325 9027
rect 17276 8996 17325 9024
rect 17276 8984 17282 8996
rect 17313 8993 17325 8996
rect 17359 8993 17371 9027
rect 17313 8987 17371 8993
rect 17773 9027 17831 9033
rect 17773 8993 17785 9027
rect 17819 9024 17831 9027
rect 17954 9024 17960 9036
rect 17819 8996 17960 9024
rect 17819 8993 17831 8996
rect 17773 8987 17831 8993
rect 17954 8984 17960 8996
rect 18012 8984 18018 9036
rect 18800 9033 18828 9064
rect 20898 9052 20904 9064
rect 20956 9052 20962 9104
rect 21468 9101 21496 9132
rect 21545 9129 21557 9163
rect 21591 9160 21603 9163
rect 22370 9160 22376 9172
rect 21591 9132 22376 9160
rect 21591 9129 21603 9132
rect 21545 9123 21603 9129
rect 22370 9120 22376 9132
rect 22428 9120 22434 9172
rect 23566 9160 23572 9172
rect 23527 9132 23572 9160
rect 23566 9120 23572 9132
rect 23624 9120 23630 9172
rect 28905 9163 28963 9169
rect 28905 9129 28917 9163
rect 28951 9160 28963 9163
rect 29086 9160 29092 9172
rect 28951 9132 29092 9160
rect 28951 9129 28963 9132
rect 28905 9123 28963 9129
rect 29086 9120 29092 9132
rect 29144 9120 29150 9172
rect 29454 9160 29460 9172
rect 29415 9132 29460 9160
rect 29454 9120 29460 9132
rect 29512 9120 29518 9172
rect 33226 9160 33232 9172
rect 31726 9132 33232 9160
rect 21453 9095 21511 9101
rect 21453 9061 21465 9095
rect 21499 9061 21511 9095
rect 30742 9092 30748 9104
rect 30703 9064 30748 9092
rect 21453 9055 21511 9061
rect 30742 9052 30748 9064
rect 30800 9052 30806 9104
rect 31726 9092 31754 9132
rect 33226 9120 33232 9132
rect 33284 9120 33290 9172
rect 31128 9064 31754 9092
rect 18785 9027 18843 9033
rect 18785 8993 18797 9027
rect 18831 8993 18843 9027
rect 18785 8987 18843 8993
rect 20717 9027 20775 9033
rect 20717 8993 20729 9027
rect 20763 9024 20775 9027
rect 20806 9024 20812 9036
rect 20763 8996 20812 9024
rect 20763 8993 20775 8996
rect 20717 8987 20775 8993
rect 19061 8959 19119 8965
rect 17144 8928 18092 8956
rect 9088 8916 9094 8928
rect 9490 8848 9496 8900
rect 9548 8888 9554 8900
rect 9585 8891 9643 8897
rect 9585 8888 9597 8891
rect 9548 8860 9597 8888
rect 9548 8848 9554 8860
rect 9585 8857 9597 8860
rect 9631 8857 9643 8891
rect 9585 8851 9643 8857
rect 18064 8888 18092 8928
rect 19061 8925 19073 8959
rect 19107 8956 19119 8959
rect 19702 8956 19708 8968
rect 19107 8928 19708 8956
rect 19107 8925 19119 8928
rect 19061 8919 19119 8925
rect 19702 8916 19708 8928
rect 19760 8916 19766 8968
rect 20732 8956 20760 8987
rect 20806 8984 20812 8996
rect 20864 8984 20870 9036
rect 22649 9027 22707 9033
rect 22649 8993 22661 9027
rect 22695 8993 22707 9027
rect 23842 9024 23848 9036
rect 23803 8996 23848 9024
rect 22649 8987 22707 8993
rect 22094 8956 22100 8968
rect 20732 8928 22100 8956
rect 22094 8916 22100 8928
rect 22152 8956 22158 8968
rect 22664 8956 22692 8987
rect 23842 8984 23848 8996
rect 23900 8984 23906 9036
rect 27062 8984 27068 9036
rect 27120 8984 27126 9036
rect 28350 8984 28356 9036
rect 28408 9024 28414 9036
rect 28721 9027 28779 9033
rect 28721 9024 28733 9027
rect 28408 8996 28733 9024
rect 28408 8984 28414 8996
rect 28721 8993 28733 8996
rect 28767 9024 28779 9027
rect 29365 9027 29423 9033
rect 29365 9024 29377 9027
rect 28767 8996 29377 9024
rect 28767 8993 28779 8996
rect 28721 8987 28779 8993
rect 29365 8993 29377 8996
rect 29411 8993 29423 9027
rect 30926 9024 30932 9036
rect 30887 8996 30932 9024
rect 29365 8987 29423 8993
rect 30926 8984 30932 8996
rect 30984 8984 30990 9036
rect 31128 9033 31156 9064
rect 32582 9052 32588 9104
rect 32640 9052 32646 9104
rect 31113 9027 31171 9033
rect 31113 8993 31125 9027
rect 31159 8993 31171 9027
rect 31113 8987 31171 8993
rect 23566 8956 23572 8968
rect 22152 8928 22692 8956
rect 23527 8928 23572 8956
rect 22152 8916 22158 8928
rect 23566 8916 23572 8928
rect 23624 8916 23630 8968
rect 25685 8959 25743 8965
rect 25685 8925 25697 8959
rect 25731 8925 25743 8959
rect 25958 8956 25964 8968
rect 25919 8928 25964 8956
rect 25685 8919 25743 8925
rect 20162 8888 20168 8900
rect 18064 8860 20168 8888
rect 3053 8823 3111 8829
rect 3053 8789 3065 8823
rect 3099 8820 3111 8823
rect 3142 8820 3148 8832
rect 3099 8792 3148 8820
rect 3099 8789 3111 8792
rect 3053 8783 3111 8789
rect 3142 8780 3148 8792
rect 3200 8780 3206 8832
rect 10686 8820 10692 8832
rect 10647 8792 10692 8820
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 18064 8829 18092 8860
rect 20162 8848 20168 8860
rect 20220 8848 20226 8900
rect 20530 8888 20536 8900
rect 20491 8860 20536 8888
rect 20530 8848 20536 8860
rect 20588 8848 20594 8900
rect 21174 8848 21180 8900
rect 21232 8888 21238 8900
rect 22833 8891 22891 8897
rect 22833 8888 22845 8891
rect 21232 8860 22845 8888
rect 21232 8848 21238 8860
rect 22833 8857 22845 8860
rect 22879 8888 22891 8891
rect 23474 8888 23480 8900
rect 22879 8860 23480 8888
rect 22879 8857 22891 8860
rect 22833 8851 22891 8857
rect 23474 8848 23480 8860
rect 23532 8888 23538 8900
rect 23753 8891 23811 8897
rect 23753 8888 23765 8891
rect 23532 8860 23765 8888
rect 23532 8848 23538 8860
rect 23753 8857 23765 8860
rect 23799 8888 23811 8891
rect 23842 8888 23848 8900
rect 23799 8860 23848 8888
rect 23799 8857 23811 8860
rect 23753 8851 23811 8857
rect 23842 8848 23848 8860
rect 23900 8848 23906 8900
rect 18049 8823 18107 8829
rect 18049 8789 18061 8823
rect 18095 8789 18107 8823
rect 18874 8820 18880 8832
rect 18835 8792 18880 8820
rect 18049 8783 18107 8789
rect 18874 8780 18880 8792
rect 18932 8780 18938 8832
rect 18966 8780 18972 8832
rect 19024 8820 19030 8832
rect 25700 8820 25728 8919
rect 25958 8916 25964 8928
rect 26016 8916 26022 8968
rect 28445 8959 28503 8965
rect 28445 8925 28457 8959
rect 28491 8956 28503 8959
rect 29086 8956 29092 8968
rect 28491 8928 29092 8956
rect 28491 8925 28503 8928
rect 28445 8919 28503 8925
rect 29086 8916 29092 8928
rect 29144 8916 29150 8968
rect 31018 8916 31024 8968
rect 31076 8956 31082 8968
rect 31573 8959 31631 8965
rect 31573 8956 31585 8959
rect 31076 8928 31585 8956
rect 31076 8916 31082 8928
rect 31573 8925 31585 8928
rect 31619 8925 31631 8959
rect 31846 8956 31852 8968
rect 31807 8928 31852 8956
rect 31573 8919 31631 8925
rect 31846 8916 31852 8928
rect 31904 8916 31910 8968
rect 32306 8916 32312 8968
rect 32364 8956 32370 8968
rect 33597 8959 33655 8965
rect 33597 8956 33609 8959
rect 32364 8928 33609 8956
rect 32364 8916 32370 8928
rect 33597 8925 33609 8928
rect 33643 8925 33655 8959
rect 33597 8919 33655 8925
rect 26050 8820 26056 8832
rect 19024 8792 19069 8820
rect 25700 8792 26056 8820
rect 19024 8780 19030 8792
rect 26050 8780 26056 8792
rect 26108 8780 26114 8832
rect 27433 8823 27491 8829
rect 27433 8789 27445 8823
rect 27479 8820 27491 8823
rect 28166 8820 28172 8832
rect 27479 8792 28172 8820
rect 27479 8789 27491 8792
rect 27433 8783 27491 8789
rect 28166 8780 28172 8792
rect 28224 8780 28230 8832
rect 28534 8820 28540 8832
rect 28495 8792 28540 8820
rect 28534 8780 28540 8792
rect 28592 8780 28598 8832
rect 1104 8730 34316 8752
rect 1104 8678 6517 8730
rect 6569 8678 6581 8730
rect 6633 8678 6645 8730
rect 6697 8678 6709 8730
rect 6761 8678 17588 8730
rect 17640 8678 17652 8730
rect 17704 8678 17716 8730
rect 17768 8678 17780 8730
rect 17832 8678 28658 8730
rect 28710 8678 28722 8730
rect 28774 8678 28786 8730
rect 28838 8678 28850 8730
rect 28902 8678 34316 8730
rect 1104 8656 34316 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 4430 8616 4436 8628
rect 4391 8588 4436 8616
rect 4430 8576 4436 8588
rect 4488 8576 4494 8628
rect 5718 8576 5724 8628
rect 5776 8616 5782 8628
rect 15933 8619 15991 8625
rect 15933 8616 15945 8619
rect 5776 8588 15945 8616
rect 5776 8576 5782 8588
rect 15933 8585 15945 8588
rect 15979 8616 15991 8619
rect 16206 8616 16212 8628
rect 15979 8588 16212 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 16301 8619 16359 8625
rect 16301 8585 16313 8619
rect 16347 8616 16359 8619
rect 16942 8616 16948 8628
rect 16347 8588 16948 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 16942 8576 16948 8588
rect 17000 8576 17006 8628
rect 17126 8576 17132 8628
rect 17184 8616 17190 8628
rect 17313 8619 17371 8625
rect 17313 8616 17325 8619
rect 17184 8588 17325 8616
rect 17184 8576 17190 8588
rect 17313 8585 17325 8588
rect 17359 8585 17371 8619
rect 17313 8579 17371 8585
rect 17954 8576 17960 8628
rect 18012 8616 18018 8628
rect 19794 8616 19800 8628
rect 18012 8588 19800 8616
rect 18012 8576 18018 8588
rect 19794 8576 19800 8588
rect 19852 8616 19858 8628
rect 20073 8619 20131 8625
rect 20073 8616 20085 8619
rect 19852 8588 20085 8616
rect 19852 8576 19858 8588
rect 20073 8585 20085 8588
rect 20119 8585 20131 8619
rect 20073 8579 20131 8585
rect 20162 8576 20168 8628
rect 20220 8616 20226 8628
rect 20220 8588 25636 8616
rect 20220 8576 20226 8588
rect 4522 8508 4528 8560
rect 4580 8548 4586 8560
rect 6822 8548 6828 8560
rect 4580 8520 6828 8548
rect 4580 8508 4586 8520
rect 6822 8508 6828 8520
rect 6880 8548 6886 8560
rect 9401 8551 9459 8557
rect 9401 8548 9413 8551
rect 6880 8520 9413 8548
rect 6880 8508 6886 8520
rect 9401 8517 9413 8520
rect 9447 8517 9459 8551
rect 11241 8551 11299 8557
rect 11241 8548 11253 8551
rect 9401 8511 9459 8517
rect 9600 8520 11253 8548
rect 3326 8480 3332 8492
rect 3287 8452 3332 8480
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 8849 8483 8907 8489
rect 8849 8449 8861 8483
rect 8895 8480 8907 8483
rect 8895 8452 9536 8480
rect 8895 8449 8907 8452
rect 8849 8443 8907 8449
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8372 1458 8424
rect 3142 8412 3148 8424
rect 3103 8384 3148 8412
rect 3142 8372 3148 8384
rect 3200 8372 3206 8424
rect 3786 8372 3792 8424
rect 3844 8412 3850 8424
rect 4249 8415 4307 8421
rect 4249 8412 4261 8415
rect 3844 8384 4261 8412
rect 3844 8372 3850 8384
rect 4249 8381 4261 8384
rect 4295 8381 4307 8415
rect 4249 8375 4307 8381
rect 8570 8344 8576 8356
rect 8531 8316 8576 8344
rect 8570 8304 8576 8316
rect 8628 8304 8634 8356
rect 9508 8344 9536 8452
rect 9600 8421 9628 8520
rect 11241 8517 11253 8520
rect 11287 8548 11299 8551
rect 11330 8548 11336 8560
rect 11287 8520 11336 8548
rect 11287 8517 11299 8520
rect 11241 8511 11299 8517
rect 11330 8508 11336 8520
rect 11388 8508 11394 8560
rect 25608 8548 25636 8588
rect 25958 8576 25964 8628
rect 26016 8616 26022 8628
rect 29733 8619 29791 8625
rect 29733 8616 29745 8619
rect 26016 8588 29745 8616
rect 26016 8576 26022 8588
rect 29733 8585 29745 8588
rect 29779 8585 29791 8619
rect 29733 8579 29791 8585
rect 31846 8576 31852 8628
rect 31904 8616 31910 8628
rect 33045 8619 33103 8625
rect 33045 8616 33057 8619
rect 31904 8588 33057 8616
rect 31904 8576 31910 8588
rect 33045 8585 33057 8588
rect 33091 8585 33103 8619
rect 33045 8579 33103 8585
rect 29089 8551 29147 8557
rect 29089 8548 29101 8551
rect 25608 8520 29101 8548
rect 29089 8517 29101 8520
rect 29135 8517 29147 8551
rect 29089 8511 29147 8517
rect 9674 8440 9680 8492
rect 9732 8480 9738 8492
rect 10597 8483 10655 8489
rect 10597 8480 10609 8483
rect 9732 8452 10609 8480
rect 9732 8440 9738 8452
rect 10597 8449 10609 8452
rect 10643 8480 10655 8483
rect 11514 8480 11520 8492
rect 10643 8452 11520 8480
rect 10643 8449 10655 8452
rect 10597 8443 10655 8449
rect 11514 8440 11520 8452
rect 11572 8480 11578 8492
rect 13173 8483 13231 8489
rect 13173 8480 13185 8483
rect 11572 8452 13185 8480
rect 11572 8440 11578 8452
rect 13173 8449 13185 8452
rect 13219 8449 13231 8483
rect 13173 8443 13231 8449
rect 20622 8440 20628 8492
rect 20680 8480 20686 8492
rect 21269 8483 21327 8489
rect 21269 8480 21281 8483
rect 20680 8452 21281 8480
rect 20680 8440 20686 8452
rect 21269 8449 21281 8452
rect 21315 8449 21327 8483
rect 30466 8480 30472 8492
rect 21269 8443 21327 8449
rect 29288 8452 30472 8480
rect 9585 8415 9643 8421
rect 9585 8381 9597 8415
rect 9631 8381 9643 8415
rect 9585 8375 9643 8381
rect 11425 8415 11483 8421
rect 11425 8381 11437 8415
rect 11471 8412 11483 8415
rect 11882 8412 11888 8424
rect 11471 8384 11888 8412
rect 11471 8381 11483 8384
rect 11425 8375 11483 8381
rect 11882 8372 11888 8384
rect 11940 8372 11946 8424
rect 15197 8415 15255 8421
rect 15197 8381 15209 8415
rect 15243 8381 15255 8415
rect 15378 8412 15384 8424
rect 15339 8384 15384 8412
rect 15197 8375 15255 8381
rect 9766 8344 9772 8356
rect 9508 8316 9772 8344
rect 9766 8304 9772 8316
rect 9824 8344 9830 8356
rect 10962 8344 10968 8356
rect 9824 8316 10968 8344
rect 9824 8304 9830 8316
rect 10962 8304 10968 8316
rect 11020 8344 11026 8356
rect 12894 8344 12900 8356
rect 11020 8316 12900 8344
rect 11020 8304 11026 8316
rect 12894 8304 12900 8316
rect 12952 8304 12958 8356
rect 15212 8344 15240 8375
rect 15378 8372 15384 8384
rect 15436 8372 15442 8424
rect 15841 8415 15899 8421
rect 15841 8381 15853 8415
rect 15887 8412 15899 8415
rect 16114 8412 16120 8424
rect 15887 8384 16120 8412
rect 15887 8381 15899 8384
rect 15841 8375 15899 8381
rect 15856 8344 15884 8375
rect 16114 8372 16120 8384
rect 16172 8372 16178 8424
rect 17034 8372 17040 8424
rect 17092 8412 17098 8424
rect 17497 8415 17555 8421
rect 17497 8412 17509 8415
rect 17092 8384 17509 8412
rect 17092 8372 17098 8384
rect 17497 8381 17509 8384
rect 17543 8381 17555 8415
rect 17954 8412 17960 8424
rect 17915 8384 17960 8412
rect 17497 8375 17555 8381
rect 17954 8372 17960 8384
rect 18012 8372 18018 8424
rect 18690 8412 18696 8424
rect 18651 8384 18696 8412
rect 18690 8372 18696 8384
rect 18748 8372 18754 8424
rect 18966 8421 18972 8424
rect 18960 8412 18972 8421
rect 18927 8384 18972 8412
rect 18960 8375 18972 8384
rect 18966 8372 18972 8375
rect 19024 8372 19030 8424
rect 20809 8415 20867 8421
rect 20809 8381 20821 8415
rect 20855 8412 20867 8415
rect 21453 8415 21511 8421
rect 21453 8412 21465 8415
rect 20855 8384 21465 8412
rect 20855 8381 20867 8384
rect 20809 8375 20867 8381
rect 21453 8381 21465 8384
rect 21499 8412 21511 8415
rect 22094 8412 22100 8424
rect 21499 8384 22100 8412
rect 21499 8381 21511 8384
rect 21453 8375 21511 8381
rect 22094 8372 22100 8384
rect 22152 8412 22158 8424
rect 22152 8384 22784 8412
rect 22152 8372 22158 8384
rect 15212 8316 15884 8344
rect 17218 8304 17224 8356
rect 17276 8344 17282 8356
rect 17865 8347 17923 8353
rect 17865 8344 17877 8347
rect 17276 8316 17877 8344
rect 17276 8304 17282 8316
rect 17865 8313 17877 8316
rect 17911 8313 17923 8347
rect 17865 8307 17923 8313
rect 18782 8304 18788 8356
rect 18840 8344 18846 8356
rect 19150 8344 19156 8356
rect 18840 8316 19156 8344
rect 18840 8304 18846 8316
rect 19150 8304 19156 8316
rect 19208 8344 19214 8356
rect 22554 8344 22560 8356
rect 19208 8316 20668 8344
rect 22515 8316 22560 8344
rect 19208 8304 19214 8316
rect 2774 8236 2780 8288
rect 2832 8276 2838 8288
rect 3234 8276 3240 8288
rect 2832 8248 2877 8276
rect 3195 8248 3240 8276
rect 2832 8236 2838 8248
rect 3234 8236 3240 8248
rect 3292 8236 3298 8288
rect 8202 8276 8208 8288
rect 8163 8248 8208 8276
rect 8202 8236 8208 8248
rect 8260 8236 8266 8288
rect 8662 8276 8668 8288
rect 8623 8248 8668 8276
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 9950 8236 9956 8288
rect 10008 8276 10014 8288
rect 10045 8279 10103 8285
rect 10045 8276 10057 8279
rect 10008 8248 10057 8276
rect 10008 8236 10014 8248
rect 10045 8245 10057 8248
rect 10091 8245 10103 8279
rect 10410 8276 10416 8288
rect 10371 8248 10416 8276
rect 10045 8239 10103 8245
rect 10410 8236 10416 8248
rect 10468 8236 10474 8288
rect 10505 8279 10563 8285
rect 10505 8245 10517 8279
rect 10551 8276 10563 8279
rect 10778 8276 10784 8288
rect 10551 8248 10784 8276
rect 10551 8245 10563 8248
rect 10505 8239 10563 8245
rect 10778 8236 10784 8248
rect 10836 8236 10842 8288
rect 12618 8276 12624 8288
rect 12579 8248 12624 8276
rect 12618 8236 12624 8248
rect 12676 8236 12682 8288
rect 12986 8276 12992 8288
rect 12947 8248 12992 8276
rect 12986 8236 12992 8248
rect 13044 8236 13050 8288
rect 13081 8279 13139 8285
rect 13081 8245 13093 8279
rect 13127 8276 13139 8279
rect 13446 8276 13452 8288
rect 13127 8248 13452 8276
rect 13127 8245 13139 8248
rect 13081 8239 13139 8245
rect 13446 8236 13452 8248
rect 13504 8236 13510 8288
rect 15381 8279 15439 8285
rect 15381 8245 15393 8279
rect 15427 8276 15439 8279
rect 15562 8276 15568 8288
rect 15427 8248 15568 8276
rect 15427 8245 15439 8248
rect 15381 8239 15439 8245
rect 15562 8236 15568 8248
rect 15620 8236 15626 8288
rect 20640 8285 20668 8316
rect 22554 8304 22560 8316
rect 22612 8304 22618 8356
rect 22756 8353 22784 8384
rect 22830 8372 22836 8424
rect 22888 8412 22894 8424
rect 23293 8415 23351 8421
rect 23293 8412 23305 8415
rect 22888 8384 23305 8412
rect 22888 8372 22894 8384
rect 23293 8381 23305 8384
rect 23339 8381 23351 8415
rect 23293 8375 23351 8381
rect 25133 8415 25191 8421
rect 25133 8381 25145 8415
rect 25179 8412 25191 8415
rect 26050 8412 26056 8424
rect 25179 8384 26056 8412
rect 25179 8381 25191 8384
rect 25133 8375 25191 8381
rect 26050 8372 26056 8384
rect 26108 8372 26114 8424
rect 28166 8412 28172 8424
rect 28127 8384 28172 8412
rect 28166 8372 28172 8384
rect 28224 8372 28230 8424
rect 29288 8421 29316 8452
rect 30466 8440 30472 8452
rect 30524 8440 30530 8492
rect 30926 8440 30932 8492
rect 30984 8480 30990 8492
rect 33226 8480 33232 8492
rect 30984 8452 31432 8480
rect 30984 8440 30990 8452
rect 31404 8424 31432 8452
rect 32048 8452 33232 8480
rect 29273 8415 29331 8421
rect 29273 8381 29285 8415
rect 29319 8381 29331 8415
rect 29273 8375 29331 8381
rect 29914 8372 29920 8424
rect 29972 8421 29978 8424
rect 29972 8415 30021 8421
rect 29972 8381 29975 8415
rect 30009 8381 30021 8415
rect 30098 8412 30104 8424
rect 30059 8384 30104 8412
rect 29972 8375 30021 8381
rect 29972 8372 29978 8375
rect 30098 8372 30104 8384
rect 30156 8372 30162 8424
rect 30190 8372 30196 8424
rect 30248 8412 30254 8424
rect 30377 8415 30435 8421
rect 30248 8384 30293 8412
rect 30248 8372 30254 8384
rect 30377 8381 30389 8415
rect 30423 8412 30435 8415
rect 31110 8412 31116 8424
rect 30423 8384 31116 8412
rect 30423 8381 30435 8384
rect 30377 8375 30435 8381
rect 31110 8372 31116 8384
rect 31168 8372 31174 8424
rect 31386 8412 31392 8424
rect 31299 8384 31392 8412
rect 31386 8372 31392 8384
rect 31444 8372 31450 8424
rect 31570 8412 31576 8424
rect 31531 8384 31576 8412
rect 31570 8372 31576 8384
rect 31628 8372 31634 8424
rect 32048 8421 32076 8452
rect 33226 8440 33232 8452
rect 33284 8440 33290 8492
rect 32033 8415 32091 8421
rect 32033 8381 32045 8415
rect 32079 8381 32091 8415
rect 33318 8412 33324 8424
rect 33279 8384 33324 8412
rect 32033 8375 32091 8381
rect 33318 8372 33324 8384
rect 33376 8372 33382 8424
rect 22741 8347 22799 8353
rect 22741 8313 22753 8347
rect 22787 8344 22799 8347
rect 22922 8344 22928 8356
rect 22787 8316 22928 8344
rect 22787 8313 22799 8316
rect 22741 8307 22799 8313
rect 22922 8304 22928 8316
rect 22980 8304 22986 8356
rect 24854 8344 24860 8356
rect 24912 8353 24918 8356
rect 24824 8316 24860 8344
rect 24854 8304 24860 8316
rect 24912 8307 24924 8353
rect 28261 8347 28319 8353
rect 28261 8313 28273 8347
rect 28307 8344 28319 8347
rect 29546 8344 29552 8356
rect 28307 8316 29552 8344
rect 28307 8313 28319 8316
rect 28261 8307 28319 8313
rect 24912 8304 24918 8307
rect 29546 8304 29552 8316
rect 29604 8304 29610 8356
rect 31478 8344 31484 8356
rect 31439 8316 31484 8344
rect 31478 8304 31484 8316
rect 31536 8304 31542 8356
rect 32950 8304 32956 8356
rect 33008 8344 33014 8356
rect 33045 8347 33103 8353
rect 33045 8344 33057 8347
rect 33008 8316 33057 8344
rect 33008 8304 33014 8316
rect 33045 8313 33057 8316
rect 33091 8313 33103 8347
rect 33045 8307 33103 8313
rect 33134 8304 33140 8356
rect 33192 8344 33198 8356
rect 33229 8347 33287 8353
rect 33229 8344 33241 8347
rect 33192 8316 33241 8344
rect 33192 8304 33198 8316
rect 33229 8313 33241 8316
rect 33275 8313 33287 8347
rect 33229 8307 33287 8313
rect 20625 8279 20683 8285
rect 20625 8245 20637 8279
rect 20671 8245 20683 8279
rect 23474 8276 23480 8288
rect 23435 8248 23480 8276
rect 20625 8239 20683 8245
rect 23474 8236 23480 8248
rect 23532 8236 23538 8288
rect 23750 8276 23756 8288
rect 23711 8248 23756 8276
rect 23750 8236 23756 8248
rect 23808 8236 23814 8288
rect 1104 8186 34316 8208
rect 1104 8134 12052 8186
rect 12104 8134 12116 8186
rect 12168 8134 12180 8186
rect 12232 8134 12244 8186
rect 12296 8134 23123 8186
rect 23175 8134 23187 8186
rect 23239 8134 23251 8186
rect 23303 8134 23315 8186
rect 23367 8134 34316 8186
rect 1104 8112 34316 8134
rect 3234 8081 3240 8084
rect 3191 8075 3240 8081
rect 3191 8041 3203 8075
rect 3237 8041 3240 8075
rect 3191 8035 3240 8041
rect 3234 8032 3240 8035
rect 3292 8032 3298 8084
rect 5350 8032 5356 8084
rect 5408 8032 5414 8084
rect 5626 8032 5632 8084
rect 5684 8072 5690 8084
rect 6319 8075 6377 8081
rect 6319 8072 6331 8075
rect 5684 8044 6331 8072
rect 5684 8032 5690 8044
rect 6319 8041 6331 8044
rect 6365 8041 6377 8075
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 6319 8035 6377 8041
rect 6932 8044 7757 8072
rect 2314 7964 2320 8016
rect 2372 7964 2378 8016
rect 5368 7990 5396 8032
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1486 7936 1492 7948
rect 1443 7908 1492 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 1486 7896 1492 7908
rect 1544 7896 1550 7948
rect 4522 7936 4528 7948
rect 4483 7908 4528 7936
rect 4522 7896 4528 7908
rect 4580 7896 4586 7948
rect 6932 7936 6960 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 7745 8035 7803 8041
rect 8113 8075 8171 8081
rect 8113 8041 8125 8075
rect 8159 8072 8171 8075
rect 8202 8072 8208 8084
rect 8159 8044 8208 8072
rect 8159 8041 8171 8044
rect 8113 8035 8171 8041
rect 8202 8032 8208 8044
rect 8260 8032 8266 8084
rect 10410 8072 10416 8084
rect 10371 8044 10416 8072
rect 10410 8032 10416 8044
rect 10468 8032 10474 8084
rect 10686 8032 10692 8084
rect 10744 8072 10750 8084
rect 10873 8075 10931 8081
rect 10873 8072 10885 8075
rect 10744 8044 10885 8072
rect 10744 8032 10750 8044
rect 10873 8041 10885 8044
rect 10919 8041 10931 8075
rect 10873 8035 10931 8041
rect 12986 8032 12992 8084
rect 13044 8072 13050 8084
rect 13081 8075 13139 8081
rect 13081 8072 13093 8075
rect 13044 8044 13093 8072
rect 13044 8032 13050 8044
rect 13081 8041 13093 8044
rect 13127 8041 13139 8075
rect 13446 8072 13452 8084
rect 13407 8044 13452 8072
rect 13081 8035 13139 8041
rect 13446 8032 13452 8044
rect 13504 8032 13510 8084
rect 16114 8072 16120 8084
rect 16075 8044 16120 8072
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 17402 8032 17408 8084
rect 17460 8072 17466 8084
rect 17681 8075 17739 8081
rect 17681 8072 17693 8075
rect 17460 8044 17693 8072
rect 17460 8032 17466 8044
rect 17681 8041 17693 8044
rect 17727 8041 17739 8075
rect 17681 8035 17739 8041
rect 18233 8075 18291 8081
rect 18233 8041 18245 8075
rect 18279 8072 18291 8075
rect 18322 8072 18328 8084
rect 18279 8044 18328 8072
rect 18279 8041 18291 8044
rect 18233 8035 18291 8041
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 24121 8075 24179 8081
rect 24121 8041 24133 8075
rect 24167 8072 24179 8075
rect 24854 8072 24860 8084
rect 24167 8044 24860 8072
rect 24167 8041 24179 8044
rect 24121 8035 24179 8041
rect 24854 8032 24860 8044
rect 24912 8032 24918 8084
rect 28534 8032 28540 8084
rect 28592 8072 28598 8084
rect 28721 8075 28779 8081
rect 28721 8072 28733 8075
rect 28592 8044 28733 8072
rect 28592 8032 28598 8044
rect 28721 8041 28733 8044
rect 28767 8041 28779 8075
rect 28721 8035 28779 8041
rect 29914 8032 29920 8084
rect 29972 8072 29978 8084
rect 30469 8075 30527 8081
rect 30469 8072 30481 8075
rect 29972 8044 30481 8072
rect 29972 8032 29978 8044
rect 30469 8041 30481 8044
rect 30515 8041 30527 8075
rect 30469 8035 30527 8041
rect 33134 8032 33140 8084
rect 33192 8072 33198 8084
rect 33505 8075 33563 8081
rect 33505 8072 33517 8075
rect 33192 8044 33517 8072
rect 33192 8032 33198 8044
rect 33505 8041 33517 8044
rect 33551 8041 33563 8075
rect 33505 8035 33563 8041
rect 9306 8004 9312 8016
rect 8128 7976 9312 8004
rect 7009 7939 7067 7945
rect 7009 7936 7021 7939
rect 6932 7908 7021 7936
rect 7009 7905 7021 7908
rect 7055 7905 7067 7939
rect 7009 7899 7067 7905
rect 7101 7939 7159 7945
rect 7101 7905 7113 7939
rect 7147 7936 7159 7939
rect 8128 7936 8156 7976
rect 9306 7964 9312 7976
rect 9364 8004 9370 8016
rect 10778 8004 10784 8016
rect 9364 7976 10088 8004
rect 10739 7976 10784 8004
rect 9364 7964 9370 7976
rect 7147 7908 8156 7936
rect 8205 7939 8263 7945
rect 7147 7905 7159 7908
rect 7101 7899 7159 7905
rect 8205 7905 8217 7939
rect 8251 7936 8263 7939
rect 8570 7936 8576 7948
rect 8251 7908 8576 7936
rect 8251 7905 8263 7908
rect 8205 7899 8263 7905
rect 8570 7896 8576 7908
rect 8628 7896 8634 7948
rect 9950 7936 9956 7948
rect 9911 7908 9956 7936
rect 9950 7896 9956 7908
rect 10008 7896 10014 7948
rect 10060 7936 10088 7976
rect 10778 7964 10784 7976
rect 10836 7964 10842 8016
rect 23293 8007 23351 8013
rect 23293 8004 23305 8007
rect 17420 7976 23305 8004
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 10060 7908 12081 7936
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7868 1823 7871
rect 2774 7868 2780 7880
rect 1811 7840 2780 7868
rect 1811 7837 1823 7840
rect 1765 7831 1823 7837
rect 2774 7828 2780 7840
rect 2832 7828 2838 7880
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7868 4951 7871
rect 5166 7868 5172 7880
rect 4939 7840 5172 7868
rect 4939 7837 4951 7840
rect 4893 7831 4951 7837
rect 5166 7828 5172 7840
rect 5224 7828 5230 7880
rect 7288 7871 7346 7877
rect 7288 7837 7300 7871
rect 7334 7837 7346 7871
rect 7288 7831 7346 7837
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7868 8447 7871
rect 8846 7868 8852 7880
rect 8435 7840 8852 7868
rect 8435 7837 8447 7840
rect 8389 7831 8447 7837
rect 7300 7800 7328 7831
rect 8846 7828 8852 7840
rect 8904 7868 8910 7880
rect 9582 7868 9588 7880
rect 8904 7840 9588 7868
rect 8904 7828 8910 7840
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 9861 7871 9919 7877
rect 9861 7837 9873 7871
rect 9907 7868 9919 7871
rect 10060 7868 10088 7908
rect 12069 7905 12081 7908
rect 12115 7905 12127 7939
rect 12069 7899 12127 7905
rect 12161 7939 12219 7945
rect 12161 7905 12173 7939
rect 12207 7936 12219 7939
rect 12618 7936 12624 7948
rect 12207 7908 12624 7936
rect 12207 7905 12219 7908
rect 12161 7899 12219 7905
rect 12618 7896 12624 7908
rect 12676 7896 12682 7948
rect 12894 7896 12900 7948
rect 12952 7936 12958 7948
rect 15004 7939 15062 7945
rect 12952 7908 13676 7936
rect 12952 7896 12958 7908
rect 10962 7868 10968 7880
rect 9907 7840 10088 7868
rect 10923 7840 10968 7868
rect 9907 7837 9919 7840
rect 9861 7831 9919 7837
rect 9692 7800 9720 7831
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 11885 7871 11943 7877
rect 11885 7837 11897 7871
rect 11931 7837 11943 7871
rect 13538 7868 13544 7880
rect 13499 7840 13544 7868
rect 11885 7831 11943 7837
rect 10134 7800 10140 7812
rect 7300 7772 10140 7800
rect 10134 7760 10140 7772
rect 10192 7800 10198 7812
rect 11900 7800 11928 7831
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 13648 7877 13676 7908
rect 15004 7905 15016 7939
rect 15050 7936 15062 7939
rect 15470 7936 15476 7948
rect 15050 7908 15476 7936
rect 15050 7905 15062 7908
rect 15004 7899 15062 7905
rect 15470 7896 15476 7908
rect 15528 7896 15534 7948
rect 17420 7945 17448 7976
rect 23293 7973 23305 7976
rect 23339 7973 23351 8007
rect 23293 7967 23351 7973
rect 28077 8007 28135 8013
rect 28077 7973 28089 8007
rect 28123 8004 28135 8007
rect 28994 8004 29000 8016
rect 28123 7976 29000 8004
rect 28123 7973 28135 7976
rect 28077 7967 28135 7973
rect 16761 7939 16819 7945
rect 16761 7905 16773 7939
rect 16807 7905 16819 7939
rect 16761 7899 16819 7905
rect 17405 7939 17463 7945
rect 17405 7905 17417 7939
rect 17451 7905 17463 7939
rect 17405 7899 17463 7905
rect 13633 7871 13691 7877
rect 13633 7837 13645 7871
rect 13679 7837 13691 7871
rect 14734 7868 14740 7880
rect 14695 7840 14740 7868
rect 13633 7831 13691 7837
rect 14734 7828 14740 7840
rect 14792 7828 14798 7880
rect 16776 7868 16804 7899
rect 18046 7896 18052 7948
rect 18104 7936 18110 7948
rect 18325 7939 18383 7945
rect 18325 7936 18337 7939
rect 18104 7908 18337 7936
rect 18104 7896 18110 7908
rect 18325 7905 18337 7908
rect 18371 7905 18383 7939
rect 18325 7899 18383 7905
rect 20346 7896 20352 7948
rect 20404 7936 20410 7948
rect 21634 7945 21640 7948
rect 20533 7939 20591 7945
rect 20533 7936 20545 7939
rect 20404 7908 20545 7936
rect 20404 7896 20410 7908
rect 20533 7905 20545 7908
rect 20579 7905 20591 7939
rect 20533 7899 20591 7905
rect 21628 7899 21640 7945
rect 21692 7936 21698 7948
rect 23385 7939 23443 7945
rect 21692 7908 21728 7936
rect 21634 7896 21640 7899
rect 21692 7896 21698 7908
rect 23385 7905 23397 7939
rect 23431 7936 23443 7939
rect 23750 7936 23756 7948
rect 23431 7908 23756 7936
rect 23431 7905 23443 7908
rect 23385 7899 23443 7905
rect 23750 7896 23756 7908
rect 23808 7896 23814 7948
rect 23845 7939 23903 7945
rect 23845 7905 23857 7939
rect 23891 7936 23903 7939
rect 26970 7936 26976 7948
rect 23891 7908 26976 7936
rect 23891 7905 23903 7908
rect 23845 7899 23903 7905
rect 26970 7896 26976 7908
rect 27028 7896 27034 7948
rect 27798 7936 27804 7948
rect 27759 7908 27804 7936
rect 27798 7896 27804 7908
rect 27856 7896 27862 7948
rect 27985 7939 28043 7945
rect 27985 7905 27997 7939
rect 28031 7936 28043 7939
rect 28166 7936 28172 7948
rect 28031 7908 28172 7936
rect 28031 7905 28043 7908
rect 27985 7899 28043 7905
rect 28166 7896 28172 7908
rect 28224 7896 28230 7948
rect 28644 7945 28672 7976
rect 28994 7964 29000 7976
rect 29052 7964 29058 8016
rect 29546 8004 29552 8016
rect 29507 7976 29552 8004
rect 29546 7964 29552 7976
rect 29604 7964 29610 8016
rect 29638 7964 29644 8016
rect 29696 8004 29702 8016
rect 29696 7976 30788 8004
rect 29696 7964 29702 7976
rect 28629 7939 28687 7945
rect 28629 7905 28641 7939
rect 28675 7905 28687 7939
rect 28629 7899 28687 7905
rect 28813 7939 28871 7945
rect 28813 7905 28825 7939
rect 28859 7936 28871 7939
rect 29270 7936 29276 7948
rect 28859 7908 29276 7936
rect 28859 7905 28871 7908
rect 28813 7899 28871 7905
rect 29270 7896 29276 7908
rect 29328 7896 29334 7948
rect 29365 7939 29423 7945
rect 29365 7905 29377 7939
rect 29411 7936 29423 7939
rect 30006 7936 30012 7948
rect 29411 7908 30012 7936
rect 29411 7905 29423 7908
rect 29365 7899 29423 7905
rect 30006 7896 30012 7908
rect 30064 7896 30070 7948
rect 30760 7945 30788 7976
rect 32876 7976 33640 8004
rect 30745 7939 30803 7945
rect 30745 7905 30757 7939
rect 30791 7905 30803 7939
rect 30745 7899 30803 7905
rect 31110 7896 31116 7948
rect 31168 7936 31174 7948
rect 31294 7936 31300 7948
rect 31168 7908 31300 7936
rect 31168 7896 31174 7908
rect 31294 7896 31300 7908
rect 31352 7896 31358 7948
rect 32306 7936 32312 7948
rect 32267 7908 32312 7936
rect 32306 7896 32312 7908
rect 32364 7896 32370 7948
rect 32876 7945 32904 7976
rect 33612 7948 33640 7976
rect 32861 7939 32919 7945
rect 32861 7905 32873 7939
rect 32907 7905 32919 7939
rect 32861 7899 32919 7905
rect 33321 7939 33379 7945
rect 33321 7905 33333 7939
rect 33367 7936 33379 7939
rect 33410 7936 33416 7948
rect 33367 7908 33416 7936
rect 33367 7905 33379 7908
rect 33321 7899 33379 7905
rect 33410 7896 33416 7908
rect 33468 7896 33474 7948
rect 33594 7896 33600 7948
rect 33652 7936 33658 7948
rect 33652 7908 33745 7936
rect 33652 7896 33658 7908
rect 17681 7871 17739 7877
rect 16776 7840 17632 7868
rect 10192 7772 11928 7800
rect 10192 7760 10198 7772
rect 16574 7760 16580 7812
rect 16632 7800 16638 7812
rect 17604 7800 17632 7840
rect 17681 7837 17693 7871
rect 17727 7868 17739 7871
rect 17954 7868 17960 7880
rect 17727 7840 17960 7868
rect 17727 7837 17739 7840
rect 17681 7831 17739 7837
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 21082 7828 21088 7880
rect 21140 7868 21146 7880
rect 21361 7871 21419 7877
rect 21361 7868 21373 7871
rect 21140 7840 21373 7868
rect 21140 7828 21146 7840
rect 21361 7837 21373 7840
rect 21407 7837 21419 7871
rect 24118 7868 24124 7880
rect 24079 7840 24124 7868
rect 21361 7831 21419 7837
rect 24118 7828 24124 7840
rect 24176 7828 24182 7880
rect 29914 7828 29920 7880
rect 29972 7868 29978 7880
rect 30653 7871 30711 7877
rect 30653 7868 30665 7871
rect 29972 7840 30665 7868
rect 29972 7828 29978 7840
rect 30653 7837 30665 7840
rect 30699 7837 30711 7871
rect 30653 7831 30711 7837
rect 31202 7828 31208 7880
rect 31260 7868 31266 7880
rect 31570 7868 31576 7880
rect 31260 7840 31576 7868
rect 31260 7828 31266 7840
rect 31570 7828 31576 7840
rect 31628 7868 31634 7880
rect 32398 7868 32404 7880
rect 31628 7840 32404 7868
rect 31628 7828 31634 7840
rect 32398 7828 32404 7840
rect 32456 7828 32462 7880
rect 16632 7772 17356 7800
rect 17604 7772 20576 7800
rect 16632 7760 16638 7772
rect 17328 7744 17356 7772
rect 7193 7735 7251 7741
rect 7193 7701 7205 7735
rect 7239 7732 7251 7735
rect 7558 7732 7564 7744
rect 7239 7704 7564 7732
rect 7239 7701 7251 7704
rect 7193 7695 7251 7701
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 9766 7732 9772 7744
rect 9727 7704 9772 7732
rect 9766 7692 9772 7704
rect 9824 7692 9830 7744
rect 11974 7732 11980 7744
rect 11935 7704 11980 7732
rect 11974 7692 11980 7704
rect 12032 7692 12038 7744
rect 16666 7732 16672 7744
rect 16627 7704 16672 7732
rect 16666 7692 16672 7704
rect 16724 7692 16730 7744
rect 17310 7732 17316 7744
rect 17223 7704 17316 7732
rect 17310 7692 17316 7704
rect 17368 7732 17374 7744
rect 17497 7735 17555 7741
rect 17497 7732 17509 7735
rect 17368 7704 17509 7732
rect 17368 7692 17374 7704
rect 17497 7701 17509 7704
rect 17543 7701 17555 7735
rect 17497 7695 17555 7701
rect 19610 7692 19616 7744
rect 19668 7732 19674 7744
rect 20441 7735 20499 7741
rect 20441 7732 20453 7735
rect 19668 7704 20453 7732
rect 19668 7692 19674 7704
rect 20441 7701 20453 7704
rect 20487 7701 20499 7735
rect 20548 7732 20576 7772
rect 23842 7760 23848 7812
rect 23900 7800 23906 7812
rect 23937 7803 23995 7809
rect 23937 7800 23949 7803
rect 23900 7772 23949 7800
rect 23900 7760 23906 7772
rect 23937 7769 23949 7772
rect 23983 7769 23995 7803
rect 23937 7763 23995 7769
rect 29549 7803 29607 7809
rect 29549 7769 29561 7803
rect 29595 7800 29607 7803
rect 30098 7800 30104 7812
rect 29595 7772 30104 7800
rect 29595 7769 29607 7772
rect 29549 7763 29607 7769
rect 30098 7760 30104 7772
rect 30156 7760 30162 7812
rect 22370 7732 22376 7744
rect 20548 7704 22376 7732
rect 20441 7695 20499 7701
rect 22370 7692 22376 7704
rect 22428 7692 22434 7744
rect 22462 7692 22468 7744
rect 22520 7732 22526 7744
rect 22741 7735 22799 7741
rect 22741 7732 22753 7735
rect 22520 7704 22753 7732
rect 22520 7692 22526 7704
rect 22741 7701 22753 7704
rect 22787 7701 22799 7735
rect 22741 7695 22799 7701
rect 33226 7692 33232 7744
rect 33284 7732 33290 7744
rect 33321 7735 33379 7741
rect 33321 7732 33333 7735
rect 33284 7704 33333 7732
rect 33284 7692 33290 7704
rect 33321 7701 33333 7704
rect 33367 7701 33379 7735
rect 33321 7695 33379 7701
rect 1104 7642 34316 7664
rect 1104 7590 6517 7642
rect 6569 7590 6581 7642
rect 6633 7590 6645 7642
rect 6697 7590 6709 7642
rect 6761 7590 17588 7642
rect 17640 7590 17652 7642
rect 17704 7590 17716 7642
rect 17768 7590 17780 7642
rect 17832 7590 28658 7642
rect 28710 7590 28722 7642
rect 28774 7590 28786 7642
rect 28838 7590 28850 7642
rect 28902 7590 34316 7642
rect 1104 7568 34316 7590
rect 5166 7528 5172 7540
rect 5127 7500 5172 7528
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 8481 7531 8539 7537
rect 8481 7497 8493 7531
rect 8527 7528 8539 7531
rect 8570 7528 8576 7540
rect 8527 7500 8576 7528
rect 8527 7497 8539 7500
rect 8481 7491 8539 7497
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 8662 7488 8668 7540
rect 8720 7528 8726 7540
rect 9033 7531 9091 7537
rect 9033 7528 9045 7531
rect 8720 7500 9045 7528
rect 8720 7488 8726 7500
rect 9033 7497 9045 7500
rect 9079 7497 9091 7531
rect 9033 7491 9091 7497
rect 15470 7488 15476 7540
rect 15528 7528 15534 7540
rect 15657 7531 15715 7537
rect 15657 7528 15669 7531
rect 15528 7500 15669 7528
rect 15528 7488 15534 7500
rect 15657 7497 15669 7500
rect 15703 7497 15715 7531
rect 19702 7528 19708 7540
rect 19663 7500 19708 7528
rect 15657 7491 15715 7497
rect 19702 7488 19708 7500
rect 19760 7488 19766 7540
rect 21174 7488 21180 7540
rect 21232 7528 21238 7540
rect 21453 7531 21511 7537
rect 21453 7528 21465 7531
rect 21232 7500 21465 7528
rect 21232 7488 21238 7500
rect 21453 7497 21465 7500
rect 21499 7497 21511 7531
rect 21453 7491 21511 7497
rect 21545 7531 21603 7537
rect 21545 7497 21557 7531
rect 21591 7528 21603 7531
rect 21634 7528 21640 7540
rect 21591 7500 21640 7528
rect 21591 7497 21603 7500
rect 21545 7491 21603 7497
rect 21634 7488 21640 7500
rect 21692 7488 21698 7540
rect 23293 7531 23351 7537
rect 23293 7497 23305 7531
rect 23339 7528 23351 7531
rect 23566 7528 23572 7540
rect 23339 7500 23572 7528
rect 23339 7497 23351 7500
rect 23293 7491 23351 7497
rect 23566 7488 23572 7500
rect 23624 7488 23630 7540
rect 24118 7528 24124 7540
rect 24079 7500 24124 7528
rect 24118 7488 24124 7500
rect 24176 7488 24182 7540
rect 28905 7531 28963 7537
rect 28905 7528 28917 7531
rect 28184 7500 28917 7528
rect 4430 7420 4436 7472
rect 4488 7460 4494 7472
rect 5442 7460 5448 7472
rect 4488 7432 5448 7460
rect 4488 7420 4494 7432
rect 5442 7420 5448 7432
rect 5500 7460 5506 7472
rect 11057 7463 11115 7469
rect 11057 7460 11069 7463
rect 5500 7432 5764 7460
rect 5500 7420 5506 7432
rect 3142 7392 3148 7404
rect 3103 7364 3148 7392
rect 3142 7352 3148 7364
rect 3200 7392 3206 7404
rect 3326 7392 3332 7404
rect 3200 7364 3332 7392
rect 3200 7352 3206 7364
rect 3326 7352 3332 7364
rect 3384 7352 3390 7404
rect 5626 7392 5632 7404
rect 5587 7364 5632 7392
rect 5626 7352 5632 7364
rect 5684 7352 5690 7404
rect 5736 7401 5764 7432
rect 10244 7432 11069 7460
rect 10244 7404 10272 7432
rect 11057 7429 11069 7432
rect 11103 7429 11115 7463
rect 11057 7423 11115 7429
rect 22370 7420 22376 7472
rect 22428 7460 22434 7472
rect 25866 7460 25872 7472
rect 22428 7432 25872 7460
rect 22428 7420 22434 7432
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 8294 7392 8300 7404
rect 7883 7364 8300 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 8294 7352 8300 7364
rect 8352 7392 8358 7404
rect 10226 7392 10232 7404
rect 8352 7364 9720 7392
rect 10187 7364 10232 7392
rect 8352 7352 8358 7364
rect 2958 7284 2964 7336
rect 3016 7324 3022 7336
rect 3053 7327 3111 7333
rect 3053 7324 3065 7327
rect 3016 7296 3065 7324
rect 3016 7284 3022 7296
rect 3053 7293 3065 7296
rect 3099 7293 3111 7327
rect 7558 7324 7564 7336
rect 7519 7296 7564 7324
rect 3053 7287 3111 7293
rect 7558 7284 7564 7296
rect 7616 7284 7622 7336
rect 8573 7327 8631 7333
rect 8573 7293 8585 7327
rect 8619 7293 8631 7327
rect 9030 7324 9036 7336
rect 8991 7296 9036 7324
rect 8573 7287 8631 7293
rect 7653 7259 7711 7265
rect 7653 7225 7665 7259
rect 7699 7256 7711 7259
rect 8588 7256 8616 7287
rect 9030 7284 9036 7296
rect 9088 7284 9094 7336
rect 9217 7327 9275 7333
rect 9217 7293 9229 7327
rect 9263 7324 9275 7327
rect 9398 7324 9404 7336
rect 9263 7296 9404 7324
rect 9263 7293 9275 7296
rect 9217 7287 9275 7293
rect 9232 7256 9260 7287
rect 9398 7284 9404 7296
rect 9456 7284 9462 7336
rect 7699 7228 9260 7256
rect 9692 7256 9720 7364
rect 10226 7352 10232 7364
rect 10284 7352 10290 7404
rect 10413 7395 10471 7401
rect 10413 7361 10425 7395
rect 10459 7392 10471 7395
rect 12621 7395 12679 7401
rect 12621 7392 12633 7395
rect 10459 7364 12633 7392
rect 10459 7361 10471 7364
rect 10413 7355 10471 7361
rect 12621 7361 12633 7364
rect 12667 7361 12679 7395
rect 12621 7355 12679 7361
rect 9766 7284 9772 7336
rect 9824 7324 9830 7336
rect 10137 7327 10195 7333
rect 10137 7324 10149 7327
rect 9824 7296 10149 7324
rect 9824 7284 9830 7296
rect 10137 7293 10149 7296
rect 10183 7293 10195 7327
rect 10137 7287 10195 7293
rect 10428 7256 10456 7355
rect 13446 7352 13452 7404
rect 13504 7392 13510 7404
rect 15562 7392 15568 7404
rect 13504 7364 14504 7392
rect 15523 7364 15568 7392
rect 13504 7352 13510 7364
rect 10778 7284 10784 7336
rect 10836 7324 10842 7336
rect 10965 7327 11023 7333
rect 10965 7324 10977 7327
rect 10836 7296 10977 7324
rect 10836 7284 10842 7296
rect 10965 7293 10977 7296
rect 11011 7293 11023 7327
rect 10965 7287 11023 7293
rect 11974 7284 11980 7336
rect 12032 7324 12038 7336
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 12032 7296 12449 7324
rect 12032 7284 12038 7296
rect 12437 7293 12449 7296
rect 12483 7293 12495 7327
rect 12437 7287 12495 7293
rect 13262 7284 13268 7336
rect 13320 7324 13326 7336
rect 13633 7327 13691 7333
rect 13633 7324 13645 7327
rect 13320 7296 13645 7324
rect 13320 7284 13326 7296
rect 13633 7293 13645 7296
rect 13679 7293 13691 7327
rect 13814 7324 13820 7336
rect 13775 7296 13820 7324
rect 13633 7287 13691 7293
rect 13814 7284 13820 7296
rect 13872 7284 13878 7336
rect 14476 7333 14504 7364
rect 15562 7352 15568 7364
rect 15620 7352 15626 7404
rect 21637 7395 21695 7401
rect 21637 7361 21649 7395
rect 21683 7392 21695 7395
rect 22649 7395 22707 7401
rect 22649 7392 22661 7395
rect 21683 7364 22661 7392
rect 21683 7361 21695 7364
rect 21637 7355 21695 7361
rect 22649 7361 22661 7364
rect 22695 7361 22707 7395
rect 22649 7355 22707 7361
rect 14461 7327 14519 7333
rect 14461 7293 14473 7327
rect 14507 7293 14519 7327
rect 15746 7324 15752 7336
rect 15707 7296 15752 7324
rect 14461 7287 14519 7293
rect 15746 7284 15752 7296
rect 15804 7284 15810 7336
rect 15841 7327 15899 7333
rect 15841 7293 15853 7327
rect 15887 7324 15899 7327
rect 16666 7324 16672 7336
rect 15887 7296 16672 7324
rect 15887 7293 15899 7296
rect 15841 7287 15899 7293
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 17126 7284 17132 7336
rect 17184 7324 17190 7336
rect 17313 7327 17371 7333
rect 17313 7324 17325 7327
rect 17184 7296 17325 7324
rect 17184 7284 17190 7296
rect 17313 7293 17325 7296
rect 17359 7293 17371 7327
rect 17313 7287 17371 7293
rect 17402 7284 17408 7336
rect 17460 7324 17466 7336
rect 17569 7327 17627 7333
rect 17569 7324 17581 7327
rect 17460 7296 17581 7324
rect 17460 7284 17466 7296
rect 17569 7293 17581 7296
rect 17615 7293 17627 7327
rect 19610 7324 19616 7336
rect 19571 7296 19616 7324
rect 17569 7287 17627 7293
rect 19610 7284 19616 7296
rect 19668 7284 19674 7336
rect 19794 7324 19800 7336
rect 19755 7296 19800 7324
rect 19794 7284 19800 7296
rect 19852 7284 19858 7336
rect 21358 7324 21364 7336
rect 21319 7296 21364 7324
rect 21358 7284 21364 7296
rect 21416 7284 21422 7336
rect 22278 7284 22284 7336
rect 22336 7324 22342 7336
rect 22557 7327 22615 7333
rect 22557 7324 22569 7327
rect 22336 7296 22569 7324
rect 22336 7284 22342 7296
rect 9692 7228 10456 7256
rect 12529 7259 12587 7265
rect 7699 7225 7711 7228
rect 7653 7219 7711 7225
rect 12529 7225 12541 7259
rect 12575 7256 12587 7259
rect 12710 7256 12716 7268
rect 12575 7228 12716 7256
rect 12575 7225 12587 7228
rect 12529 7219 12587 7225
rect 12710 7216 12716 7228
rect 12768 7256 12774 7268
rect 14553 7259 14611 7265
rect 14553 7256 14565 7259
rect 12768 7228 14565 7256
rect 12768 7216 12774 7228
rect 14553 7225 14565 7228
rect 14599 7225 14611 7259
rect 14553 7219 14611 7225
rect 1854 7148 1860 7200
rect 1912 7188 1918 7200
rect 2593 7191 2651 7197
rect 2593 7188 2605 7191
rect 1912 7160 2605 7188
rect 1912 7148 1918 7160
rect 2593 7157 2605 7160
rect 2639 7157 2651 7191
rect 2593 7151 2651 7157
rect 2961 7191 3019 7197
rect 2961 7157 2973 7191
rect 3007 7188 3019 7191
rect 3234 7188 3240 7200
rect 3007 7160 3240 7188
rect 3007 7157 3019 7160
rect 2961 7151 3019 7157
rect 3234 7148 3240 7160
rect 3292 7148 3298 7200
rect 5534 7188 5540 7200
rect 5495 7160 5540 7188
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 7190 7188 7196 7200
rect 7151 7160 7196 7188
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 9582 7148 9588 7200
rect 9640 7188 9646 7200
rect 9769 7191 9827 7197
rect 9769 7188 9781 7191
rect 9640 7160 9781 7188
rect 9640 7148 9646 7160
rect 9769 7157 9781 7160
rect 9815 7157 9827 7191
rect 9769 7151 9827 7157
rect 11790 7148 11796 7200
rect 11848 7188 11854 7200
rect 12069 7191 12127 7197
rect 12069 7188 12081 7191
rect 11848 7160 12081 7188
rect 11848 7148 11854 7160
rect 12069 7157 12081 7160
rect 12115 7157 12127 7191
rect 13998 7188 14004 7200
rect 13959 7160 14004 7188
rect 12069 7151 12127 7157
rect 13998 7148 14004 7160
rect 14056 7148 14062 7200
rect 18046 7148 18052 7200
rect 18104 7188 18110 7200
rect 18693 7191 18751 7197
rect 18693 7188 18705 7191
rect 18104 7160 18705 7188
rect 18104 7148 18110 7160
rect 18693 7157 18705 7160
rect 18739 7157 18751 7191
rect 22388 7188 22416 7296
rect 22557 7293 22569 7296
rect 22603 7293 22615 7327
rect 22557 7287 22615 7293
rect 22741 7327 22799 7333
rect 22741 7293 22753 7327
rect 22787 7293 22799 7327
rect 22741 7287 22799 7293
rect 22462 7216 22468 7268
rect 22520 7256 22526 7268
rect 22756 7256 22784 7287
rect 22922 7284 22928 7336
rect 22980 7324 22986 7336
rect 23400 7333 23428 7432
rect 25866 7420 25872 7432
rect 25924 7420 25930 7472
rect 23474 7352 23480 7404
rect 23532 7392 23538 7404
rect 23532 7364 24716 7392
rect 23532 7352 23538 7364
rect 23201 7327 23259 7333
rect 23201 7324 23213 7327
rect 22980 7296 23213 7324
rect 22980 7284 22986 7296
rect 23201 7293 23213 7296
rect 23247 7293 23259 7327
rect 23201 7287 23259 7293
rect 23385 7327 23443 7333
rect 23385 7293 23397 7327
rect 23431 7293 23443 7327
rect 23385 7287 23443 7293
rect 23750 7284 23756 7336
rect 23808 7324 23814 7336
rect 24688 7333 24716 7364
rect 24029 7327 24087 7333
rect 24029 7324 24041 7327
rect 23808 7296 24041 7324
rect 23808 7284 23814 7296
rect 24029 7293 24041 7296
rect 24075 7293 24087 7327
rect 24029 7287 24087 7293
rect 24213 7327 24271 7333
rect 24213 7293 24225 7327
rect 24259 7293 24271 7327
rect 24213 7287 24271 7293
rect 24673 7327 24731 7333
rect 24673 7293 24685 7327
rect 24719 7293 24731 7327
rect 24673 7287 24731 7293
rect 27985 7327 28043 7333
rect 27985 7293 27997 7327
rect 28031 7324 28043 7327
rect 28074 7324 28080 7336
rect 28031 7296 28080 7324
rect 28031 7293 28043 7296
rect 27985 7287 28043 7293
rect 22520 7228 22784 7256
rect 22520 7216 22526 7228
rect 22922 7188 22928 7200
rect 22388 7160 22928 7188
rect 18693 7151 18751 7157
rect 22922 7148 22928 7160
rect 22980 7188 22986 7200
rect 24228 7188 24256 7287
rect 28074 7284 28080 7296
rect 28132 7284 28138 7336
rect 28184 7333 28212 7500
rect 28905 7497 28917 7500
rect 28951 7497 28963 7531
rect 29914 7528 29920 7540
rect 29875 7500 29920 7528
rect 28905 7491 28963 7497
rect 29914 7488 29920 7500
rect 29972 7488 29978 7540
rect 32398 7488 32404 7540
rect 32456 7528 32462 7540
rect 33229 7531 33287 7537
rect 33229 7528 33241 7531
rect 32456 7500 33241 7528
rect 32456 7488 32462 7500
rect 33229 7497 33241 7500
rect 33275 7497 33287 7531
rect 33229 7491 33287 7497
rect 28534 7420 28540 7472
rect 28592 7460 28598 7472
rect 28997 7463 29055 7469
rect 28997 7460 29009 7463
rect 28592 7432 29009 7460
rect 28592 7420 28598 7432
rect 28997 7429 29009 7432
rect 29043 7429 29055 7463
rect 28997 7423 29055 7429
rect 29822 7420 29828 7472
rect 29880 7420 29886 7472
rect 30006 7420 30012 7472
rect 30064 7460 30070 7472
rect 33410 7460 33416 7472
rect 30064 7432 33416 7460
rect 30064 7420 30070 7432
rect 33410 7420 33416 7432
rect 33468 7420 33474 7472
rect 28905 7395 28963 7401
rect 28905 7361 28917 7395
rect 28951 7392 28963 7395
rect 29840 7392 29868 7420
rect 28951 7364 29868 7392
rect 28951 7361 28963 7364
rect 28905 7355 28963 7361
rect 30466 7352 30472 7404
rect 30524 7392 30530 7404
rect 30653 7395 30711 7401
rect 30653 7392 30665 7395
rect 30524 7364 30665 7392
rect 30524 7352 30530 7364
rect 30653 7361 30665 7364
rect 30699 7392 30711 7395
rect 31110 7392 31116 7404
rect 30699 7364 31116 7392
rect 30699 7361 30711 7364
rect 30653 7355 30711 7361
rect 31110 7352 31116 7364
rect 31168 7352 31174 7404
rect 28169 7327 28227 7333
rect 28169 7293 28181 7327
rect 28215 7293 28227 7327
rect 28169 7287 28227 7293
rect 28261 7327 28319 7333
rect 28261 7293 28273 7327
rect 28307 7324 28319 7327
rect 28442 7324 28448 7336
rect 28307 7296 28448 7324
rect 28307 7293 28319 7296
rect 28261 7287 28319 7293
rect 28442 7284 28448 7296
rect 28500 7284 28506 7336
rect 29086 7324 29092 7336
rect 29047 7296 29092 7324
rect 29086 7284 29092 7296
rect 29144 7284 29150 7336
rect 29546 7284 29552 7336
rect 29604 7324 29610 7336
rect 29825 7327 29883 7333
rect 29825 7324 29837 7327
rect 29604 7296 29837 7324
rect 29604 7284 29610 7296
rect 29825 7293 29837 7296
rect 29871 7293 29883 7327
rect 29825 7287 29883 7293
rect 30009 7327 30067 7333
rect 30009 7293 30021 7327
rect 30055 7293 30067 7327
rect 30558 7324 30564 7336
rect 30519 7296 30564 7324
rect 30009 7287 30067 7293
rect 28718 7256 28724 7268
rect 28679 7228 28724 7256
rect 28718 7216 28724 7228
rect 28776 7216 28782 7268
rect 29730 7216 29736 7268
rect 29788 7256 29794 7268
rect 30024 7256 30052 7287
rect 30558 7284 30564 7296
rect 30616 7284 30622 7336
rect 31202 7324 31208 7336
rect 31163 7296 31208 7324
rect 31202 7284 31208 7296
rect 31260 7284 31266 7336
rect 31294 7284 31300 7336
rect 31352 7324 31358 7336
rect 31352 7296 31397 7324
rect 31352 7284 31358 7296
rect 33318 7265 33324 7268
rect 29788 7228 30052 7256
rect 33045 7259 33103 7265
rect 29788 7216 29794 7228
rect 33045 7225 33057 7259
rect 33091 7225 33103 7259
rect 33045 7219 33103 7225
rect 33261 7259 33324 7265
rect 33261 7225 33273 7259
rect 33307 7225 33324 7259
rect 33261 7219 33324 7225
rect 22980 7160 24256 7188
rect 24857 7191 24915 7197
rect 22980 7148 22986 7160
rect 24857 7157 24869 7191
rect 24903 7188 24915 7191
rect 26050 7188 26056 7200
rect 24903 7160 26056 7188
rect 24903 7157 24915 7160
rect 24857 7151 24915 7157
rect 26050 7148 26056 7160
rect 26108 7148 26114 7200
rect 26234 7148 26240 7200
rect 26292 7188 26298 7200
rect 27801 7191 27859 7197
rect 27801 7188 27813 7191
rect 26292 7160 27813 7188
rect 26292 7148 26298 7160
rect 27801 7157 27813 7160
rect 27847 7157 27859 7191
rect 27801 7151 27859 7157
rect 31386 7148 31392 7200
rect 31444 7188 31450 7200
rect 33060 7188 33088 7219
rect 33318 7216 33324 7219
rect 33376 7216 33382 7268
rect 31444 7160 33088 7188
rect 31444 7148 31450 7160
rect 1104 7098 34316 7120
rect 1104 7046 12052 7098
rect 12104 7046 12116 7098
rect 12168 7046 12180 7098
rect 12232 7046 12244 7098
rect 12296 7046 23123 7098
rect 23175 7046 23187 7098
rect 23239 7046 23251 7098
rect 23303 7046 23315 7098
rect 23367 7046 34316 7098
rect 1104 7024 34316 7046
rect 2314 6944 2320 6996
rect 2372 6984 2378 6996
rect 2682 6984 2688 6996
rect 2372 6956 2688 6984
rect 2372 6944 2378 6956
rect 2682 6944 2688 6956
rect 2740 6944 2746 6996
rect 10689 6987 10747 6993
rect 10689 6953 10701 6987
rect 10735 6984 10747 6987
rect 10778 6984 10784 6996
rect 10735 6956 10784 6984
rect 10735 6953 10747 6956
rect 10689 6947 10747 6953
rect 10778 6944 10784 6956
rect 10836 6944 10842 6996
rect 12805 6987 12863 6993
rect 12805 6953 12817 6987
rect 12851 6984 12863 6987
rect 13538 6984 13544 6996
rect 12851 6956 13544 6984
rect 12851 6953 12863 6956
rect 12805 6947 12863 6953
rect 13538 6944 13544 6956
rect 13596 6944 13602 6996
rect 17865 6987 17923 6993
rect 17865 6953 17877 6987
rect 17911 6984 17923 6987
rect 17954 6984 17960 6996
rect 17911 6956 17960 6984
rect 17911 6953 17923 6956
rect 17865 6947 17923 6953
rect 17954 6944 17960 6956
rect 18012 6944 18018 6996
rect 27893 6987 27951 6993
rect 27893 6953 27905 6987
rect 27939 6984 27951 6987
rect 28718 6984 28724 6996
rect 27939 6956 28724 6984
rect 27939 6953 27951 6956
rect 27893 6947 27951 6953
rect 28718 6944 28724 6956
rect 28776 6944 28782 6996
rect 33594 6984 33600 6996
rect 33555 6956 33600 6984
rect 33594 6944 33600 6956
rect 33652 6944 33658 6996
rect 2332 6902 2360 6944
rect 5261 6919 5319 6925
rect 5261 6885 5273 6919
rect 5307 6916 5319 6919
rect 5626 6916 5632 6928
rect 5307 6888 5632 6916
rect 5307 6885 5319 6888
rect 5261 6879 5319 6885
rect 5626 6876 5632 6888
rect 5684 6876 5690 6928
rect 10594 6876 10600 6928
rect 10652 6916 10658 6928
rect 11057 6919 11115 6925
rect 11057 6916 11069 6919
rect 10652 6888 11069 6916
rect 10652 6876 10658 6888
rect 11057 6885 11069 6888
rect 11103 6885 11115 6919
rect 11057 6879 11115 6885
rect 13262 6876 13268 6928
rect 13320 6916 13326 6928
rect 13725 6919 13783 6925
rect 13725 6916 13737 6919
rect 13320 6888 13737 6916
rect 13320 6876 13326 6888
rect 13725 6885 13737 6888
rect 13771 6885 13783 6919
rect 13725 6879 13783 6885
rect 17126 6876 17132 6928
rect 17184 6916 17190 6928
rect 18690 6916 18696 6928
rect 17184 6888 18696 6916
rect 17184 6876 17190 6888
rect 18690 6876 18696 6888
rect 18748 6916 18754 6928
rect 19518 6916 19524 6928
rect 18748 6888 19524 6916
rect 18748 6876 18754 6888
rect 19518 6876 19524 6888
rect 19576 6876 19582 6928
rect 25958 6916 25964 6928
rect 25608 6888 25964 6916
rect 1854 6848 1860 6860
rect 1815 6820 1860 6848
rect 1854 6808 1860 6820
rect 1912 6808 1918 6860
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6848 5411 6851
rect 5534 6848 5540 6860
rect 5399 6820 5540 6848
rect 5399 6817 5411 6820
rect 5353 6811 5411 6817
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 11330 6808 11336 6860
rect 11388 6848 11394 6860
rect 11977 6851 12035 6857
rect 11977 6848 11989 6851
rect 11388 6820 11989 6848
rect 11388 6808 11394 6820
rect 11977 6817 11989 6820
rect 12023 6817 12035 6851
rect 12710 6848 12716 6860
rect 12671 6820 12716 6848
rect 11977 6811 12035 6817
rect 12710 6808 12716 6820
rect 12768 6808 12774 6860
rect 12897 6851 12955 6857
rect 12897 6817 12909 6851
rect 12943 6817 12955 6851
rect 12897 6811 12955 6817
rect 1394 6740 1400 6792
rect 1452 6780 1458 6792
rect 1489 6783 1547 6789
rect 1489 6780 1501 6783
rect 1452 6752 1501 6780
rect 1452 6740 1458 6752
rect 1489 6749 1501 6752
rect 1535 6780 1547 6783
rect 5442 6780 5448 6792
rect 1535 6752 2728 6780
rect 5403 6752 5448 6780
rect 1535 6749 1547 6752
rect 1489 6743 1547 6749
rect 2700 6712 2728 6752
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 10962 6740 10968 6792
rect 11020 6780 11026 6792
rect 11149 6783 11207 6789
rect 11149 6780 11161 6783
rect 11020 6752 11161 6780
rect 11020 6740 11026 6752
rect 11149 6749 11161 6752
rect 11195 6749 11207 6783
rect 11149 6743 11207 6749
rect 11241 6783 11299 6789
rect 11241 6749 11253 6783
rect 11287 6749 11299 6783
rect 11241 6743 11299 6749
rect 4522 6712 4528 6724
rect 2700 6684 4528 6712
rect 4522 6672 4528 6684
rect 4580 6672 4586 6724
rect 10042 6672 10048 6724
rect 10100 6712 10106 6724
rect 11256 6712 11284 6743
rect 11606 6740 11612 6792
rect 11664 6780 11670 6792
rect 12912 6780 12940 6811
rect 13170 6808 13176 6860
rect 13228 6848 13234 6860
rect 13357 6851 13415 6857
rect 13357 6848 13369 6851
rect 13228 6820 13369 6848
rect 13228 6808 13234 6820
rect 13357 6817 13369 6820
rect 13403 6817 13415 6851
rect 13357 6811 13415 6817
rect 13541 6851 13599 6857
rect 13541 6817 13553 6851
rect 13587 6848 13599 6851
rect 13630 6848 13636 6860
rect 13587 6820 13636 6848
rect 13587 6817 13599 6820
rect 13541 6811 13599 6817
rect 13630 6808 13636 6820
rect 13688 6808 13694 6860
rect 15749 6851 15807 6857
rect 15749 6817 15761 6851
rect 15795 6848 15807 6851
rect 15930 6848 15936 6860
rect 15795 6820 15936 6848
rect 15795 6817 15807 6820
rect 15749 6811 15807 6817
rect 15930 6808 15936 6820
rect 15988 6808 15994 6860
rect 16206 6808 16212 6860
rect 16264 6848 16270 6860
rect 16669 6851 16727 6857
rect 16669 6848 16681 6851
rect 16264 6820 16681 6848
rect 16264 6808 16270 6820
rect 16669 6817 16681 6820
rect 16715 6817 16727 6851
rect 16669 6811 16727 6817
rect 16758 6808 16764 6860
rect 16816 6848 16822 6860
rect 17865 6851 17923 6857
rect 17865 6848 17877 6851
rect 16816 6820 16861 6848
rect 17788 6820 17877 6848
rect 16816 6808 16822 6820
rect 11664 6752 12940 6780
rect 15473 6783 15531 6789
rect 11664 6740 11670 6752
rect 15473 6749 15485 6783
rect 15519 6780 15531 6783
rect 16482 6780 16488 6792
rect 15519 6752 16488 6780
rect 15519 6749 15531 6752
rect 15473 6743 15531 6749
rect 16482 6740 16488 6752
rect 16540 6740 16546 6792
rect 13354 6712 13360 6724
rect 10100 6684 13360 6712
rect 10100 6672 10106 6684
rect 13354 6672 13360 6684
rect 13412 6712 13418 6724
rect 13538 6712 13544 6724
rect 13412 6684 13544 6712
rect 13412 6672 13418 6684
rect 13538 6672 13544 6684
rect 13596 6672 13602 6724
rect 15378 6672 15384 6724
rect 15436 6712 15442 6724
rect 17788 6712 17816 6820
rect 17865 6817 17877 6820
rect 17911 6817 17923 6851
rect 18046 6848 18052 6860
rect 18007 6820 18052 6848
rect 17865 6811 17923 6817
rect 18046 6808 18052 6820
rect 18104 6808 18110 6860
rect 19058 6848 19064 6860
rect 19019 6820 19064 6848
rect 19058 6808 19064 6820
rect 19116 6808 19122 6860
rect 20625 6851 20683 6857
rect 20625 6817 20637 6851
rect 20671 6848 20683 6851
rect 21177 6851 21235 6857
rect 21177 6848 21189 6851
rect 20671 6820 21189 6848
rect 20671 6817 20683 6820
rect 20625 6811 20683 6817
rect 21177 6817 21189 6820
rect 21223 6817 21235 6851
rect 21177 6811 21235 6817
rect 21266 6808 21272 6860
rect 21324 6848 21330 6860
rect 21913 6851 21971 6857
rect 21324 6820 21369 6848
rect 21324 6808 21330 6820
rect 21913 6817 21925 6851
rect 21959 6848 21971 6851
rect 23474 6848 23480 6860
rect 21959 6820 23480 6848
rect 21959 6817 21971 6820
rect 21913 6811 21971 6817
rect 23474 6808 23480 6820
rect 23532 6808 23538 6860
rect 23753 6851 23811 6857
rect 23753 6817 23765 6851
rect 23799 6848 23811 6851
rect 23934 6848 23940 6860
rect 23799 6820 23940 6848
rect 23799 6817 23811 6820
rect 23753 6811 23811 6817
rect 23934 6808 23940 6820
rect 23992 6808 23998 6860
rect 25608 6857 25636 6888
rect 25958 6876 25964 6888
rect 26016 6876 26022 6928
rect 32582 6876 32588 6928
rect 32640 6876 32646 6928
rect 25593 6851 25651 6857
rect 25593 6817 25605 6851
rect 25639 6817 25651 6851
rect 25593 6811 25651 6817
rect 26970 6808 26976 6860
rect 27028 6808 27034 6860
rect 27798 6848 27804 6860
rect 27356 6820 27804 6848
rect 18785 6783 18843 6789
rect 18785 6749 18797 6783
rect 18831 6780 18843 6783
rect 20070 6780 20076 6792
rect 18831 6752 20076 6780
rect 18831 6749 18843 6752
rect 18785 6743 18843 6749
rect 20070 6740 20076 6752
rect 20128 6740 20134 6792
rect 20346 6780 20352 6792
rect 20307 6752 20352 6780
rect 20346 6740 20352 6752
rect 20404 6740 20410 6792
rect 23842 6780 23848 6792
rect 23803 6752 23848 6780
rect 23842 6740 23848 6752
rect 23900 6740 23906 6792
rect 24026 6780 24032 6792
rect 23987 6752 24032 6780
rect 24026 6740 24032 6752
rect 24084 6740 24090 6792
rect 25869 6783 25927 6789
rect 25869 6749 25881 6783
rect 25915 6780 25927 6783
rect 26234 6780 26240 6792
rect 25915 6752 26240 6780
rect 25915 6749 25927 6752
rect 25869 6743 25927 6749
rect 26234 6740 26240 6752
rect 26292 6740 26298 6792
rect 27356 6789 27384 6820
rect 27798 6808 27804 6820
rect 27856 6808 27862 6860
rect 28721 6851 28779 6857
rect 28721 6817 28733 6851
rect 28767 6817 28779 6851
rect 28721 6811 28779 6817
rect 28905 6851 28963 6857
rect 28905 6817 28917 6851
rect 28951 6848 28963 6851
rect 29270 6848 29276 6860
rect 28951 6820 29276 6848
rect 28951 6817 28963 6820
rect 28905 6811 28963 6817
rect 27341 6783 27399 6789
rect 27341 6749 27353 6783
rect 27387 6749 27399 6783
rect 28736 6780 28764 6811
rect 29270 6808 29276 6820
rect 29328 6808 29334 6860
rect 29362 6808 29368 6860
rect 29420 6848 29426 6860
rect 29549 6851 29607 6857
rect 29420 6820 29465 6848
rect 29420 6808 29426 6820
rect 29549 6817 29561 6851
rect 29595 6848 29607 6851
rect 30006 6848 30012 6860
rect 29595 6820 30012 6848
rect 29595 6817 29607 6820
rect 29549 6811 29607 6817
rect 30006 6808 30012 6820
rect 30064 6808 30070 6860
rect 29457 6783 29515 6789
rect 29457 6780 29469 6783
rect 28736 6752 29469 6780
rect 27341 6743 27399 6749
rect 29457 6749 29469 6752
rect 29503 6749 29515 6783
rect 29457 6743 29515 6749
rect 31018 6740 31024 6792
rect 31076 6780 31082 6792
rect 31570 6780 31576 6792
rect 31076 6752 31576 6780
rect 31076 6740 31082 6752
rect 31570 6740 31576 6752
rect 31628 6780 31634 6792
rect 31849 6783 31907 6789
rect 31849 6780 31861 6783
rect 31628 6752 31861 6780
rect 31628 6740 31634 6752
rect 31849 6749 31861 6752
rect 31895 6749 31907 6783
rect 31849 6743 31907 6749
rect 32125 6783 32183 6789
rect 32125 6749 32137 6783
rect 32171 6780 32183 6783
rect 33134 6780 33140 6792
rect 32171 6752 33140 6780
rect 32171 6749 32183 6752
rect 32125 6743 32183 6749
rect 33134 6740 33140 6752
rect 33192 6740 33198 6792
rect 19610 6712 19616 6724
rect 15436 6684 19616 6712
rect 15436 6672 15442 6684
rect 19610 6672 19616 6684
rect 19668 6672 19674 6724
rect 20533 6715 20591 6721
rect 20533 6712 20545 6715
rect 19720 6684 20545 6712
rect 2958 6604 2964 6656
rect 3016 6644 3022 6656
rect 3283 6647 3341 6653
rect 3283 6644 3295 6647
rect 3016 6616 3295 6644
rect 3016 6604 3022 6616
rect 3283 6613 3295 6616
rect 3329 6613 3341 6647
rect 3283 6607 3341 6613
rect 4246 6604 4252 6656
rect 4304 6644 4310 6656
rect 4893 6647 4951 6653
rect 4893 6644 4905 6647
rect 4304 6616 4905 6644
rect 4304 6604 4310 6616
rect 4893 6613 4905 6616
rect 4939 6613 4951 6647
rect 4893 6607 4951 6613
rect 12161 6647 12219 6653
rect 12161 6613 12173 6647
rect 12207 6644 12219 6647
rect 12342 6644 12348 6656
rect 12207 6616 12348 6644
rect 12207 6613 12219 6616
rect 12161 6607 12219 6613
rect 12342 6604 12348 6616
rect 12400 6604 12406 6656
rect 15562 6644 15568 6656
rect 15523 6616 15568 6644
rect 15562 6604 15568 6616
rect 15620 6604 15626 6656
rect 15657 6647 15715 6653
rect 15657 6613 15669 6647
rect 15703 6644 15715 6647
rect 15746 6644 15752 6656
rect 15703 6616 15752 6644
rect 15703 6613 15715 6616
rect 15657 6607 15715 6613
rect 15746 6604 15752 6616
rect 15804 6644 15810 6656
rect 18690 6644 18696 6656
rect 15804 6616 18696 6644
rect 15804 6604 15810 6616
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 18874 6644 18880 6656
rect 18835 6616 18880 6644
rect 18874 6604 18880 6616
rect 18932 6604 18938 6656
rect 18966 6604 18972 6656
rect 19024 6644 19030 6656
rect 19720 6644 19748 6684
rect 20533 6681 20545 6684
rect 20579 6712 20591 6715
rect 22554 6712 22560 6724
rect 20579 6684 22560 6712
rect 20579 6681 20591 6684
rect 20533 6675 20591 6681
rect 22554 6672 22560 6684
rect 22612 6672 22618 6724
rect 19024 6616 19748 6644
rect 19024 6604 19030 6616
rect 20254 6604 20260 6656
rect 20312 6644 20318 6656
rect 20441 6647 20499 6653
rect 20441 6644 20453 6647
rect 20312 6616 20453 6644
rect 20312 6604 20318 6616
rect 20441 6613 20453 6616
rect 20487 6613 20499 6647
rect 21726 6644 21732 6656
rect 21687 6616 21732 6644
rect 20441 6607 20499 6613
rect 21726 6604 21732 6616
rect 21784 6604 21790 6656
rect 23937 6647 23995 6653
rect 23937 6613 23949 6647
rect 23983 6644 23995 6647
rect 24394 6644 24400 6656
rect 23983 6616 24400 6644
rect 23983 6613 23995 6616
rect 23937 6607 23995 6613
rect 24394 6604 24400 6616
rect 24452 6604 24458 6656
rect 28258 6604 28264 6656
rect 28316 6644 28322 6656
rect 28813 6647 28871 6653
rect 28813 6644 28825 6647
rect 28316 6616 28825 6644
rect 28316 6604 28322 6616
rect 28813 6613 28825 6616
rect 28859 6613 28871 6647
rect 28813 6607 28871 6613
rect 1104 6554 34316 6576
rect 1104 6502 6517 6554
rect 6569 6502 6581 6554
rect 6633 6502 6645 6554
rect 6697 6502 6709 6554
rect 6761 6502 17588 6554
rect 17640 6502 17652 6554
rect 17704 6502 17716 6554
rect 17768 6502 17780 6554
rect 17832 6502 28658 6554
rect 28710 6502 28722 6554
rect 28774 6502 28786 6554
rect 28838 6502 28850 6554
rect 28902 6502 34316 6554
rect 1104 6480 34316 6502
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 5675 6443 5733 6449
rect 5675 6440 5687 6443
rect 5592 6412 5687 6440
rect 5592 6400 5598 6412
rect 5675 6409 5687 6412
rect 5721 6409 5733 6443
rect 9398 6440 9404 6452
rect 9359 6412 9404 6440
rect 5675 6403 5733 6409
rect 9398 6400 9404 6412
rect 9456 6400 9462 6452
rect 10962 6440 10968 6452
rect 10923 6412 10968 6440
rect 10962 6400 10968 6412
rect 11020 6400 11026 6452
rect 13170 6440 13176 6452
rect 12636 6412 13176 6440
rect 4246 6304 4252 6316
rect 4207 6276 4252 6304
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 4522 6304 4528 6316
rect 4356 6276 4528 6304
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 4356 6236 4384 6276
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 6914 6304 6920 6316
rect 6875 6276 6920 6304
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 7190 6304 7196 6316
rect 7151 6276 7196 6304
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 10042 6304 10048 6316
rect 10003 6276 10048 6304
rect 10042 6264 10048 6276
rect 10100 6264 10106 6316
rect 12636 6248 12664 6412
rect 13170 6400 13176 6412
rect 13228 6400 13234 6452
rect 13357 6443 13415 6449
rect 13357 6409 13369 6443
rect 13403 6440 13415 6443
rect 13446 6440 13452 6452
rect 13403 6412 13452 6440
rect 13403 6409 13415 6412
rect 13357 6403 13415 6409
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 13538 6400 13544 6452
rect 13596 6440 13602 6452
rect 16206 6440 16212 6452
rect 13596 6412 13952 6440
rect 16167 6412 16212 6440
rect 13596 6400 13602 6412
rect 12802 6372 12808 6384
rect 12715 6344 12808 6372
rect 12802 6332 12808 6344
rect 12860 6372 12866 6384
rect 13722 6372 13728 6384
rect 12860 6344 13728 6372
rect 12860 6332 12866 6344
rect 13722 6332 13728 6344
rect 13780 6332 13786 6384
rect 13630 6304 13636 6316
rect 12912 6276 13636 6304
rect 3927 6208 4384 6236
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 8202 6196 8208 6248
rect 8260 6236 8266 6248
rect 8260 6208 9996 6236
rect 8260 6196 8266 6208
rect 5258 6128 5264 6180
rect 5316 6128 5322 6180
rect 8941 6171 8999 6177
rect 8941 6137 8953 6171
rect 8987 6168 8999 6171
rect 9490 6168 9496 6180
rect 8987 6140 9496 6168
rect 8987 6137 8999 6140
rect 8941 6131 8999 6137
rect 9490 6128 9496 6140
rect 9548 6168 9554 6180
rect 9861 6171 9919 6177
rect 9861 6168 9873 6171
rect 9548 6140 9873 6168
rect 9548 6128 9554 6140
rect 9861 6137 9873 6140
rect 9907 6137 9919 6171
rect 9968 6168 9996 6208
rect 10226 6196 10232 6248
rect 10284 6236 10290 6248
rect 10873 6239 10931 6245
rect 10873 6236 10885 6239
rect 10284 6208 10885 6236
rect 10284 6196 10290 6208
rect 10873 6205 10885 6208
rect 10919 6205 10931 6239
rect 12618 6236 12624 6248
rect 12531 6208 12624 6236
rect 10873 6199 10931 6205
rect 12618 6196 12624 6208
rect 12676 6236 12682 6248
rect 12912 6245 12940 6276
rect 13630 6264 13636 6276
rect 13688 6304 13694 6316
rect 13924 6313 13952 6412
rect 16206 6400 16212 6412
rect 16264 6400 16270 6452
rect 21082 6440 21088 6452
rect 19996 6412 21088 6440
rect 13817 6307 13875 6313
rect 13817 6304 13829 6307
rect 13688 6276 13829 6304
rect 13688 6264 13694 6276
rect 13817 6273 13829 6276
rect 13863 6273 13875 6307
rect 13817 6267 13875 6273
rect 13909 6307 13967 6313
rect 13909 6273 13921 6307
rect 13955 6273 13967 6307
rect 13909 6267 13967 6273
rect 14734 6264 14740 6316
rect 14792 6304 14798 6316
rect 14829 6307 14887 6313
rect 14829 6304 14841 6307
rect 14792 6276 14841 6304
rect 14792 6264 14798 6276
rect 14829 6273 14841 6276
rect 14875 6273 14887 6307
rect 19518 6304 19524 6316
rect 19479 6276 19524 6304
rect 14829 6267 14887 6273
rect 19518 6264 19524 6276
rect 19576 6304 19582 6316
rect 19996 6313 20024 6412
rect 21082 6400 21088 6412
rect 21140 6440 21146 6452
rect 21726 6440 21732 6452
rect 21140 6412 21732 6440
rect 21140 6400 21146 6412
rect 21726 6400 21732 6412
rect 21784 6400 21790 6452
rect 22554 6400 22560 6452
rect 22612 6440 22618 6452
rect 22741 6443 22799 6449
rect 22741 6440 22753 6443
rect 22612 6412 22753 6440
rect 22612 6400 22618 6412
rect 22741 6409 22753 6412
rect 22787 6409 22799 6443
rect 29270 6440 29276 6452
rect 29231 6412 29276 6440
rect 22741 6403 22799 6409
rect 29270 6400 29276 6412
rect 29328 6400 29334 6452
rect 29362 6400 29368 6452
rect 29420 6440 29426 6452
rect 30009 6443 30067 6449
rect 30009 6440 30021 6443
rect 29420 6412 30021 6440
rect 29420 6400 29426 6412
rect 30009 6409 30021 6412
rect 30055 6409 30067 6443
rect 30009 6403 30067 6409
rect 30193 6443 30251 6449
rect 30193 6409 30205 6443
rect 30239 6440 30251 6443
rect 30558 6440 30564 6452
rect 30239 6412 30564 6440
rect 30239 6409 30251 6412
rect 30193 6403 30251 6409
rect 30558 6400 30564 6412
rect 30616 6400 30622 6452
rect 33134 6400 33140 6452
rect 33192 6440 33198 6452
rect 33229 6443 33287 6449
rect 33229 6440 33241 6443
rect 33192 6412 33241 6440
rect 33192 6400 33198 6412
rect 33229 6409 33241 6412
rect 33275 6409 33287 6443
rect 33229 6403 33287 6409
rect 19981 6307 20039 6313
rect 19981 6304 19993 6307
rect 19576 6276 19993 6304
rect 19576 6264 19582 6276
rect 19981 6273 19993 6276
rect 20027 6273 20039 6307
rect 19981 6267 20039 6273
rect 22557 6307 22615 6313
rect 22557 6273 22569 6307
rect 22603 6304 22615 6307
rect 23014 6304 23020 6316
rect 22603 6276 23020 6304
rect 22603 6273 22615 6276
rect 22557 6267 22615 6273
rect 23014 6264 23020 6276
rect 23072 6264 23078 6316
rect 23658 6264 23664 6316
rect 23716 6304 23722 6316
rect 29181 6307 29239 6313
rect 23716 6276 23888 6304
rect 23716 6264 23722 6276
rect 12713 6239 12771 6245
rect 12713 6236 12725 6239
rect 12676 6208 12725 6236
rect 12676 6196 12682 6208
rect 12713 6205 12725 6208
rect 12759 6205 12771 6239
rect 12713 6199 12771 6205
rect 12897 6239 12955 6245
rect 12897 6205 12909 6239
rect 12943 6205 12955 6239
rect 12897 6199 12955 6205
rect 13725 6239 13783 6245
rect 13725 6205 13737 6239
rect 13771 6236 13783 6239
rect 13998 6236 14004 6248
rect 13771 6208 14004 6236
rect 13771 6205 13783 6208
rect 13725 6199 13783 6205
rect 13998 6196 14004 6208
rect 14056 6196 14062 6248
rect 15096 6239 15154 6245
rect 15096 6205 15108 6239
rect 15142 6236 15154 6239
rect 15562 6236 15568 6248
rect 15142 6208 15568 6236
rect 15142 6205 15154 6208
rect 15096 6199 15154 6205
rect 15562 6196 15568 6208
rect 15620 6196 15626 6248
rect 18874 6196 18880 6248
rect 18932 6236 18938 6248
rect 20254 6245 20260 6248
rect 19254 6239 19312 6245
rect 19254 6236 19266 6239
rect 18932 6208 19266 6236
rect 18932 6196 18938 6208
rect 19254 6205 19266 6208
rect 19300 6205 19312 6239
rect 20248 6236 20260 6245
rect 20215 6208 20260 6236
rect 19254 6199 19312 6205
rect 20248 6199 20260 6208
rect 20254 6196 20260 6199
rect 20312 6196 20318 6248
rect 23860 6245 23888 6276
rect 29181 6273 29193 6307
rect 29227 6304 29239 6307
rect 29270 6304 29276 6316
rect 29227 6276 29276 6304
rect 29227 6273 29239 6276
rect 29181 6267 29239 6273
rect 29270 6264 29276 6276
rect 29328 6304 29334 6316
rect 29328 6276 30880 6304
rect 29328 6264 29334 6276
rect 22833 6239 22891 6245
rect 22833 6205 22845 6239
rect 22879 6236 22891 6239
rect 23753 6239 23811 6245
rect 23753 6236 23765 6239
rect 22879 6208 23765 6236
rect 22879 6205 22891 6208
rect 22833 6199 22891 6205
rect 23753 6205 23765 6208
rect 23799 6205 23811 6239
rect 23753 6199 23811 6205
rect 23845 6239 23903 6245
rect 23845 6205 23857 6239
rect 23891 6205 23903 6239
rect 23845 6199 23903 6205
rect 24305 6239 24363 6245
rect 24305 6205 24317 6239
rect 24351 6205 24363 6239
rect 24305 6199 24363 6205
rect 13078 6168 13084 6180
rect 9968 6140 13084 6168
rect 9861 6131 9919 6137
rect 13078 6128 13084 6140
rect 13136 6128 13142 6180
rect 16114 6128 16120 6180
rect 16172 6168 16178 6180
rect 22462 6168 22468 6180
rect 16172 6140 22468 6168
rect 16172 6128 16178 6140
rect 22462 6128 22468 6140
rect 22520 6128 22526 6180
rect 24320 6168 24348 6199
rect 24394 6196 24400 6248
rect 24452 6236 24458 6248
rect 24561 6239 24619 6245
rect 24561 6236 24573 6239
rect 24452 6208 24573 6236
rect 24452 6196 24458 6208
rect 24561 6205 24573 6208
rect 24607 6205 24619 6239
rect 28074 6236 28080 6248
rect 28035 6208 28080 6236
rect 24561 6199 24619 6205
rect 28074 6196 28080 6208
rect 28132 6196 28138 6248
rect 28258 6236 28264 6248
rect 28219 6208 28264 6236
rect 28258 6196 28264 6208
rect 28316 6196 28322 6248
rect 28353 6239 28411 6245
rect 28353 6205 28365 6239
rect 28399 6236 28411 6239
rect 28442 6236 28448 6248
rect 28399 6208 28448 6236
rect 28399 6205 28411 6208
rect 28353 6199 28411 6205
rect 28442 6196 28448 6208
rect 28500 6196 28506 6248
rect 29365 6239 29423 6245
rect 29365 6205 29377 6239
rect 29411 6205 29423 6239
rect 29365 6199 29423 6205
rect 29457 6239 29515 6245
rect 29457 6205 29469 6239
rect 29503 6236 29515 6239
rect 30466 6236 30472 6248
rect 29503 6208 30472 6236
rect 29503 6205 29515 6208
rect 29457 6199 29515 6205
rect 26050 6168 26056 6180
rect 24320 6140 26056 6168
rect 26050 6128 26056 6140
rect 26108 6128 26114 6180
rect 29380 6168 29408 6199
rect 30466 6196 30472 6208
rect 30524 6196 30530 6248
rect 30852 6245 30880 6276
rect 30837 6239 30895 6245
rect 30837 6205 30849 6239
rect 30883 6205 30895 6239
rect 30837 6199 30895 6205
rect 31481 6239 31539 6245
rect 31481 6205 31493 6239
rect 31527 6236 31539 6239
rect 31662 6236 31668 6248
rect 31527 6208 31668 6236
rect 31527 6205 31539 6208
rect 31481 6199 31539 6205
rect 31662 6196 31668 6208
rect 31720 6196 31726 6248
rect 32950 6196 32956 6248
rect 33008 6236 33014 6248
rect 33045 6239 33103 6245
rect 33045 6236 33057 6239
rect 33008 6208 33057 6236
rect 33008 6196 33014 6208
rect 33045 6205 33057 6208
rect 33091 6205 33103 6239
rect 33226 6236 33232 6248
rect 33187 6208 33232 6236
rect 33045 6199 33103 6205
rect 33226 6196 33232 6208
rect 33284 6196 33290 6248
rect 29638 6168 29644 6180
rect 29380 6140 29644 6168
rect 29638 6128 29644 6140
rect 29696 6128 29702 6180
rect 29730 6128 29736 6180
rect 29788 6168 29794 6180
rect 30161 6171 30219 6177
rect 30161 6168 30173 6171
rect 29788 6140 30173 6168
rect 29788 6128 29794 6140
rect 30161 6137 30173 6140
rect 30207 6168 30219 6171
rect 30377 6171 30435 6177
rect 30207 6137 30236 6168
rect 30161 6131 30236 6137
rect 30377 6137 30389 6171
rect 30423 6168 30435 6171
rect 31294 6168 31300 6180
rect 30423 6140 31300 6168
rect 30423 6137 30435 6140
rect 30377 6131 30435 6137
rect 9766 6100 9772 6112
rect 9727 6072 9772 6100
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 18141 6103 18199 6109
rect 18141 6069 18153 6103
rect 18187 6100 18199 6103
rect 18414 6100 18420 6112
rect 18187 6072 18420 6100
rect 18187 6069 18199 6072
rect 18141 6063 18199 6069
rect 18414 6060 18420 6072
rect 18472 6060 18478 6112
rect 21358 6100 21364 6112
rect 21319 6072 21364 6100
rect 21358 6060 21364 6072
rect 21416 6060 21422 6112
rect 22554 6100 22560 6112
rect 22515 6072 22560 6100
rect 22554 6060 22560 6072
rect 22612 6060 22618 6112
rect 25685 6103 25743 6109
rect 25685 6069 25697 6103
rect 25731 6100 25743 6103
rect 25958 6100 25964 6112
rect 25731 6072 25964 6100
rect 25731 6069 25743 6072
rect 25685 6063 25743 6069
rect 25958 6060 25964 6072
rect 26016 6060 26022 6112
rect 27798 6060 27804 6112
rect 27856 6100 27862 6112
rect 27893 6103 27951 6109
rect 27893 6100 27905 6103
rect 27856 6072 27905 6100
rect 27856 6060 27862 6072
rect 27893 6069 27905 6072
rect 27939 6069 27951 6103
rect 30208 6100 30236 6131
rect 31294 6128 31300 6140
rect 31352 6128 31358 6180
rect 30929 6103 30987 6109
rect 30929 6100 30941 6103
rect 30208 6072 30941 6100
rect 27893 6063 27951 6069
rect 30929 6069 30941 6072
rect 30975 6069 30987 6103
rect 30929 6063 30987 6069
rect 31573 6103 31631 6109
rect 31573 6069 31585 6103
rect 31619 6100 31631 6103
rect 31662 6100 31668 6112
rect 31619 6072 31668 6100
rect 31619 6069 31631 6072
rect 31573 6063 31631 6069
rect 31662 6060 31668 6072
rect 31720 6060 31726 6112
rect 1104 6010 34316 6032
rect 1104 5958 12052 6010
rect 12104 5958 12116 6010
rect 12168 5958 12180 6010
rect 12232 5958 12244 6010
rect 12296 5958 23123 6010
rect 23175 5958 23187 6010
rect 23239 5958 23251 6010
rect 23303 5958 23315 6010
rect 23367 5958 34316 6010
rect 1104 5936 34316 5958
rect 2958 5896 2964 5908
rect 2919 5868 2964 5896
rect 2958 5856 2964 5868
rect 3016 5856 3022 5908
rect 5626 5856 5632 5908
rect 5684 5905 5690 5908
rect 5684 5899 5733 5905
rect 5684 5865 5687 5899
rect 5721 5865 5733 5899
rect 5684 5859 5733 5865
rect 8205 5899 8263 5905
rect 8205 5865 8217 5899
rect 8251 5896 8263 5899
rect 9766 5896 9772 5908
rect 8251 5868 9772 5896
rect 8251 5865 8263 5868
rect 8205 5859 8263 5865
rect 5684 5856 5690 5859
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 10505 5899 10563 5905
rect 10505 5865 10517 5899
rect 10551 5896 10563 5899
rect 12618 5896 12624 5908
rect 10551 5868 12624 5896
rect 10551 5865 10563 5868
rect 10505 5859 10563 5865
rect 5258 5788 5264 5840
rect 5316 5828 5322 5840
rect 8389 5831 8447 5837
rect 5316 5800 6118 5828
rect 5316 5788 5322 5800
rect 8389 5797 8401 5831
rect 8435 5828 8447 5831
rect 10520 5828 10548 5859
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 15930 5896 15936 5908
rect 15891 5868 15936 5896
rect 15930 5856 15936 5868
rect 15988 5856 15994 5908
rect 16482 5896 16488 5908
rect 16443 5868 16488 5896
rect 16482 5856 16488 5868
rect 16540 5856 16546 5908
rect 20070 5896 20076 5908
rect 20031 5868 20076 5896
rect 20070 5856 20076 5868
rect 20128 5856 20134 5908
rect 20346 5856 20352 5908
rect 20404 5896 20410 5908
rect 20625 5899 20683 5905
rect 20625 5896 20637 5899
rect 20404 5868 20637 5896
rect 20404 5856 20410 5868
rect 20625 5865 20637 5868
rect 20671 5865 20683 5899
rect 26970 5896 26976 5908
rect 20625 5859 20683 5865
rect 26804 5868 26976 5896
rect 11790 5828 11796 5840
rect 8435 5800 10548 5828
rect 11751 5800 11796 5828
rect 8435 5797 8447 5800
rect 8389 5791 8447 5797
rect 11790 5788 11796 5800
rect 11848 5788 11854 5840
rect 13078 5828 13084 5840
rect 12991 5800 13084 5828
rect 13078 5788 13084 5800
rect 13136 5828 13142 5840
rect 13722 5828 13728 5840
rect 13136 5800 13728 5828
rect 13136 5788 13142 5800
rect 13722 5788 13728 5800
rect 13780 5788 13786 5840
rect 16206 5788 16212 5840
rect 16264 5828 16270 5840
rect 22186 5828 22192 5840
rect 16264 5800 16712 5828
rect 16264 5788 16270 5800
rect 8570 5760 8576 5772
rect 8531 5732 8576 5760
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 9490 5720 9496 5772
rect 9548 5760 9554 5772
rect 9769 5763 9827 5769
rect 9769 5760 9781 5763
rect 9548 5732 9781 5760
rect 9548 5720 9554 5732
rect 9769 5729 9781 5732
rect 9815 5729 9827 5763
rect 9769 5723 9827 5729
rect 10137 5763 10195 5769
rect 10137 5729 10149 5763
rect 10183 5760 10195 5763
rect 10226 5760 10232 5772
rect 10183 5732 10232 5760
rect 10183 5729 10195 5732
rect 10137 5723 10195 5729
rect 10226 5720 10232 5732
rect 10284 5720 10290 5772
rect 10410 5760 10416 5772
rect 10371 5732 10416 5760
rect 10410 5720 10416 5732
rect 10468 5720 10474 5772
rect 16025 5763 16083 5769
rect 16025 5729 16037 5763
rect 16071 5760 16083 5763
rect 16114 5760 16120 5772
rect 16071 5732 16120 5760
rect 16071 5729 16083 5732
rect 16025 5723 16083 5729
rect 16114 5720 16120 5732
rect 16172 5720 16178 5772
rect 16684 5769 16712 5800
rect 17328 5800 22192 5828
rect 17328 5769 17356 5800
rect 22186 5788 22192 5800
rect 22244 5788 22250 5840
rect 22364 5831 22422 5837
rect 22364 5797 22376 5831
rect 22410 5828 22422 5831
rect 22554 5828 22560 5840
rect 22410 5800 22560 5828
rect 22410 5797 22422 5800
rect 22364 5791 22422 5797
rect 22554 5788 22560 5800
rect 22612 5788 22618 5840
rect 26804 5814 26832 5868
rect 26970 5856 26976 5868
rect 27028 5896 27034 5908
rect 27522 5896 27528 5908
rect 27028 5868 27528 5896
rect 27028 5856 27034 5868
rect 27522 5856 27528 5868
rect 27580 5896 27586 5908
rect 29270 5896 29276 5908
rect 27580 5868 28304 5896
rect 29231 5868 29276 5896
rect 27580 5856 27586 5868
rect 27798 5828 27804 5840
rect 27759 5800 27804 5828
rect 27798 5788 27804 5800
rect 27856 5788 27862 5840
rect 28276 5814 28304 5868
rect 29270 5856 29276 5868
rect 29328 5856 29334 5908
rect 30374 5788 30380 5840
rect 30432 5828 30438 5840
rect 30929 5831 30987 5837
rect 30929 5828 30941 5831
rect 30432 5800 30941 5828
rect 30432 5788 30438 5800
rect 30929 5797 30941 5800
rect 30975 5828 30987 5831
rect 31478 5828 31484 5840
rect 30975 5800 31484 5828
rect 30975 5797 30987 5800
rect 30929 5791 30987 5797
rect 31478 5788 31484 5800
rect 31536 5788 31542 5840
rect 32858 5788 32864 5840
rect 32916 5788 32922 5840
rect 16485 5763 16543 5769
rect 16485 5729 16497 5763
rect 16531 5729 16543 5763
rect 16485 5723 16543 5729
rect 16669 5763 16727 5769
rect 16669 5729 16681 5763
rect 16715 5729 16727 5763
rect 16669 5723 16727 5729
rect 17313 5763 17371 5769
rect 17313 5729 17325 5763
rect 17359 5729 17371 5763
rect 17313 5723 17371 5729
rect 3050 5692 3056 5704
rect 3011 5664 3056 5692
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 3234 5692 3240 5704
rect 3195 5664 3240 5692
rect 3234 5652 3240 5664
rect 3292 5652 3298 5704
rect 7098 5692 7104 5704
rect 7059 5664 7104 5692
rect 7098 5652 7104 5664
rect 7156 5652 7162 5704
rect 7469 5695 7527 5701
rect 7469 5661 7481 5695
rect 7515 5692 7527 5695
rect 9306 5692 9312 5704
rect 7515 5664 9312 5692
rect 7515 5661 7527 5664
rect 7469 5655 7527 5661
rect 9306 5652 9312 5664
rect 9364 5692 9370 5704
rect 11517 5695 11575 5701
rect 11517 5692 11529 5695
rect 9364 5664 11529 5692
rect 9364 5652 9370 5664
rect 11517 5661 11529 5664
rect 11563 5692 11575 5695
rect 12342 5692 12348 5704
rect 11563 5664 12348 5692
rect 11563 5661 11575 5664
rect 11517 5655 11575 5661
rect 12342 5652 12348 5664
rect 12400 5692 12406 5704
rect 14734 5692 14740 5704
rect 12400 5664 14740 5692
rect 12400 5652 12406 5664
rect 14734 5652 14740 5664
rect 14792 5652 14798 5704
rect 15378 5652 15384 5704
rect 15436 5692 15442 5704
rect 16500 5692 16528 5723
rect 17402 5720 17408 5772
rect 17460 5760 17466 5772
rect 17460 5732 17505 5760
rect 17460 5720 17466 5732
rect 17954 5720 17960 5772
rect 18012 5760 18018 5772
rect 18233 5763 18291 5769
rect 18233 5760 18245 5763
rect 18012 5732 18245 5760
rect 18012 5720 18018 5732
rect 18233 5729 18245 5732
rect 18279 5729 18291 5763
rect 18233 5723 18291 5729
rect 18414 5720 18420 5772
rect 18472 5760 18478 5772
rect 19981 5763 20039 5769
rect 19981 5760 19993 5763
rect 18472 5732 19993 5760
rect 18472 5720 18478 5732
rect 19981 5729 19993 5732
rect 20027 5729 20039 5763
rect 19981 5723 20039 5729
rect 20165 5763 20223 5769
rect 20165 5729 20177 5763
rect 20211 5760 20223 5763
rect 20625 5763 20683 5769
rect 20625 5760 20637 5763
rect 20211 5732 20637 5760
rect 20211 5729 20223 5732
rect 20165 5723 20223 5729
rect 20625 5729 20637 5732
rect 20671 5729 20683 5763
rect 20625 5723 20683 5729
rect 20809 5763 20867 5769
rect 20809 5729 20821 5763
rect 20855 5760 20867 5763
rect 21358 5760 21364 5772
rect 20855 5732 21364 5760
rect 20855 5729 20867 5732
rect 20809 5723 20867 5729
rect 17589 5695 17647 5701
rect 17589 5692 17601 5695
rect 15436 5664 16528 5692
rect 17328 5664 17601 5692
rect 15436 5652 15442 5664
rect 17328 5636 17356 5664
rect 17589 5661 17601 5664
rect 17635 5661 17647 5695
rect 17589 5655 17647 5661
rect 19610 5652 19616 5704
rect 19668 5692 19674 5704
rect 20180 5692 20208 5723
rect 21358 5720 21364 5732
rect 21416 5720 21422 5772
rect 24121 5763 24179 5769
rect 24121 5729 24133 5763
rect 24167 5760 24179 5763
rect 24302 5760 24308 5772
rect 24167 5732 24308 5760
rect 24167 5729 24179 5732
rect 24121 5723 24179 5729
rect 24302 5720 24308 5732
rect 24360 5720 24366 5772
rect 19668 5664 20208 5692
rect 22097 5695 22155 5701
rect 19668 5652 19674 5664
rect 22097 5661 22109 5695
rect 22143 5661 22155 5695
rect 22097 5655 22155 5661
rect 25317 5695 25375 5701
rect 25317 5661 25329 5695
rect 25363 5661 25375 5695
rect 25590 5692 25596 5704
rect 25551 5664 25596 5692
rect 25317 5655 25375 5661
rect 17310 5584 17316 5636
rect 17368 5584 17374 5636
rect 17494 5624 17500 5636
rect 17455 5596 17500 5624
rect 17494 5584 17500 5596
rect 17552 5584 17558 5636
rect 21726 5584 21732 5636
rect 21784 5624 21790 5636
rect 22112 5624 22140 5655
rect 24029 5627 24087 5633
rect 24029 5624 24041 5627
rect 21784 5596 22140 5624
rect 23032 5596 24041 5624
rect 21784 5584 21790 5596
rect 2590 5556 2596 5568
rect 2551 5528 2596 5556
rect 2590 5516 2596 5528
rect 2648 5516 2654 5568
rect 13265 5559 13323 5565
rect 13265 5525 13277 5559
rect 13311 5556 13323 5559
rect 13354 5556 13360 5568
rect 13311 5528 13360 5556
rect 13311 5525 13323 5528
rect 13265 5519 13323 5525
rect 13354 5516 13360 5528
rect 13412 5516 13418 5568
rect 18138 5556 18144 5568
rect 18099 5528 18144 5556
rect 18138 5516 18144 5528
rect 18196 5516 18202 5568
rect 19058 5516 19064 5568
rect 19116 5556 19122 5568
rect 23032 5556 23060 5596
rect 24029 5593 24041 5596
rect 24075 5593 24087 5627
rect 24029 5587 24087 5593
rect 23474 5556 23480 5568
rect 19116 5528 23060 5556
rect 23435 5528 23480 5556
rect 19116 5516 19122 5528
rect 23474 5516 23480 5528
rect 23532 5516 23538 5568
rect 25332 5556 25360 5655
rect 25590 5652 25596 5664
rect 25648 5652 25654 5704
rect 26050 5652 26056 5704
rect 26108 5692 26114 5704
rect 27525 5695 27583 5701
rect 27525 5692 27537 5695
rect 26108 5664 27537 5692
rect 26108 5652 26114 5664
rect 27525 5661 27537 5664
rect 27571 5692 27583 5695
rect 31570 5692 31576 5704
rect 27571 5664 31576 5692
rect 27571 5661 27583 5664
rect 27525 5655 27583 5661
rect 31570 5652 31576 5664
rect 31628 5692 31634 5704
rect 31849 5695 31907 5701
rect 31849 5692 31861 5695
rect 31628 5664 31861 5692
rect 31628 5652 31634 5664
rect 31849 5661 31861 5664
rect 31895 5661 31907 5695
rect 32122 5692 32128 5704
rect 32083 5664 32128 5692
rect 31849 5655 31907 5661
rect 32122 5652 32128 5664
rect 32180 5652 32186 5704
rect 26050 5556 26056 5568
rect 25332 5528 26056 5556
rect 26050 5516 26056 5528
rect 26108 5516 26114 5568
rect 27062 5556 27068 5568
rect 27023 5528 27068 5556
rect 27062 5516 27068 5528
rect 27120 5516 27126 5568
rect 29086 5516 29092 5568
rect 29144 5556 29150 5568
rect 31021 5559 31079 5565
rect 31021 5556 31033 5559
rect 29144 5528 31033 5556
rect 29144 5516 29150 5528
rect 31021 5525 31033 5528
rect 31067 5525 31079 5559
rect 31021 5519 31079 5525
rect 32306 5516 32312 5568
rect 32364 5556 32370 5568
rect 33597 5559 33655 5565
rect 33597 5556 33609 5559
rect 32364 5528 33609 5556
rect 32364 5516 32370 5528
rect 33597 5525 33609 5528
rect 33643 5525 33655 5559
rect 33597 5519 33655 5525
rect 1104 5466 34316 5488
rect 1104 5414 6517 5466
rect 6569 5414 6581 5466
rect 6633 5414 6645 5466
rect 6697 5414 6709 5466
rect 6761 5414 17588 5466
rect 17640 5414 17652 5466
rect 17704 5414 17716 5466
rect 17768 5414 17780 5466
rect 17832 5414 28658 5466
rect 28710 5414 28722 5466
rect 28774 5414 28786 5466
rect 28838 5414 28850 5466
rect 28902 5414 34316 5466
rect 1104 5392 34316 5414
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 3191 5355 3249 5361
rect 3191 5352 3203 5355
rect 3108 5324 3203 5352
rect 3108 5312 3114 5324
rect 3191 5321 3203 5324
rect 3237 5321 3249 5355
rect 3191 5315 3249 5321
rect 5905 5355 5963 5361
rect 5905 5321 5917 5355
rect 5951 5352 5963 5355
rect 7098 5352 7104 5364
rect 5951 5324 7104 5352
rect 5951 5321 5963 5324
rect 5905 5315 5963 5321
rect 7098 5312 7104 5324
rect 7156 5312 7162 5364
rect 8570 5312 8576 5364
rect 8628 5352 8634 5364
rect 9125 5355 9183 5361
rect 9125 5352 9137 5355
rect 8628 5324 9137 5352
rect 8628 5312 8634 5324
rect 9125 5321 9137 5324
rect 9171 5321 9183 5355
rect 10594 5352 10600 5364
rect 10555 5324 10600 5352
rect 9125 5315 9183 5321
rect 10594 5312 10600 5324
rect 10652 5312 10658 5364
rect 13449 5355 13507 5361
rect 13449 5321 13461 5355
rect 13495 5352 13507 5355
rect 13630 5352 13636 5364
rect 13495 5324 13636 5352
rect 13495 5321 13507 5324
rect 13449 5315 13507 5321
rect 13630 5312 13636 5324
rect 13688 5312 13694 5364
rect 20530 5312 20536 5364
rect 20588 5352 20594 5364
rect 20717 5355 20775 5361
rect 20717 5352 20729 5355
rect 20588 5324 20729 5352
rect 20588 5312 20594 5324
rect 20717 5321 20729 5324
rect 20763 5321 20775 5355
rect 20717 5315 20775 5321
rect 22186 5312 22192 5364
rect 22244 5352 22250 5364
rect 22649 5355 22707 5361
rect 22649 5352 22661 5355
rect 22244 5324 22661 5352
rect 22244 5312 22250 5324
rect 22649 5321 22661 5324
rect 22695 5321 22707 5355
rect 22649 5315 22707 5321
rect 23014 5312 23020 5364
rect 23072 5352 23078 5364
rect 23293 5355 23351 5361
rect 23293 5352 23305 5355
rect 23072 5324 23305 5352
rect 23072 5312 23078 5324
rect 23293 5321 23305 5324
rect 23339 5321 23351 5355
rect 23293 5315 23351 5321
rect 24026 5312 24032 5364
rect 24084 5352 24090 5364
rect 24213 5355 24271 5361
rect 24213 5352 24225 5355
rect 24084 5324 24225 5352
rect 24084 5312 24090 5324
rect 24213 5321 24225 5324
rect 24259 5321 24271 5355
rect 24213 5315 24271 5321
rect 25501 5355 25559 5361
rect 25501 5321 25513 5355
rect 25547 5352 25559 5355
rect 25590 5352 25596 5364
rect 25547 5324 25596 5352
rect 25547 5321 25559 5324
rect 25501 5315 25559 5321
rect 25590 5312 25596 5324
rect 25648 5312 25654 5364
rect 31941 5355 31999 5361
rect 31941 5321 31953 5355
rect 31987 5352 31999 5355
rect 32122 5352 32128 5364
rect 31987 5324 32128 5352
rect 31987 5321 31999 5324
rect 31941 5315 31999 5321
rect 32122 5312 32128 5324
rect 32180 5312 32186 5364
rect 25682 5244 25688 5296
rect 25740 5284 25746 5296
rect 30929 5287 30987 5293
rect 25740 5256 26096 5284
rect 25740 5244 25746 5256
rect 1394 5216 1400 5228
rect 1355 5188 1400 5216
rect 1394 5176 1400 5188
rect 1452 5176 1458 5228
rect 1765 5219 1823 5225
rect 1765 5185 1777 5219
rect 1811 5216 1823 5219
rect 2590 5216 2596 5228
rect 1811 5188 2596 5216
rect 1811 5185 1823 5188
rect 1765 5179 1823 5185
rect 2590 5176 2596 5188
rect 2648 5176 2654 5228
rect 5350 5216 5356 5228
rect 5311 5188 5356 5216
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 5445 5219 5503 5225
rect 5445 5185 5457 5219
rect 5491 5216 5503 5219
rect 5626 5216 5632 5228
rect 5491 5188 5632 5216
rect 5491 5185 5503 5188
rect 5445 5179 5503 5185
rect 5626 5176 5632 5188
rect 5684 5176 5690 5228
rect 9493 5219 9551 5225
rect 9493 5185 9505 5219
rect 9539 5216 9551 5219
rect 10318 5216 10324 5228
rect 9539 5188 10324 5216
rect 9539 5185 9551 5188
rect 9493 5179 9551 5185
rect 10318 5176 10324 5188
rect 10376 5176 10382 5228
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5216 16175 5219
rect 16298 5216 16304 5228
rect 16163 5188 16304 5216
rect 16163 5185 16175 5188
rect 16117 5179 16175 5185
rect 16298 5176 16304 5188
rect 16356 5176 16362 5228
rect 17126 5176 17132 5228
rect 17184 5216 17190 5228
rect 17313 5219 17371 5225
rect 17313 5216 17325 5219
rect 17184 5188 17325 5216
rect 17184 5176 17190 5188
rect 17313 5185 17325 5188
rect 17359 5185 17371 5219
rect 17313 5179 17371 5185
rect 20806 5176 20812 5228
rect 20864 5216 20870 5228
rect 20901 5219 20959 5225
rect 20901 5216 20913 5219
rect 20864 5188 20913 5216
rect 20864 5176 20870 5188
rect 20901 5185 20913 5188
rect 20947 5185 20959 5219
rect 25958 5216 25964 5228
rect 20901 5179 20959 5185
rect 23216 5188 24164 5216
rect 25919 5188 25964 5216
rect 2682 5108 2688 5160
rect 2740 5148 2746 5160
rect 9309 5151 9367 5157
rect 2740 5120 2820 5148
rect 2740 5108 2746 5120
rect 2792 5080 2820 5120
rect 9309 5117 9321 5151
rect 9355 5148 9367 5151
rect 9398 5148 9404 5160
rect 9355 5120 9404 5148
rect 9355 5117 9367 5120
rect 9309 5111 9367 5117
rect 9398 5108 9404 5120
rect 9456 5108 9462 5160
rect 9585 5151 9643 5157
rect 9585 5117 9597 5151
rect 9631 5148 9643 5151
rect 10229 5151 10287 5157
rect 10229 5148 10241 5151
rect 9631 5120 10241 5148
rect 9631 5117 9643 5120
rect 9585 5111 9643 5117
rect 10229 5117 10241 5120
rect 10275 5148 10287 5151
rect 10410 5148 10416 5160
rect 10275 5120 10416 5148
rect 10275 5117 10287 5120
rect 10229 5111 10287 5117
rect 5166 5080 5172 5092
rect 2792 5066 5172 5080
rect 2806 5052 5172 5066
rect 5166 5040 5172 5052
rect 5224 5040 5230 5092
rect 9214 5040 9220 5092
rect 9272 5080 9278 5092
rect 9600 5080 9628 5111
rect 10410 5108 10416 5120
rect 10468 5108 10474 5160
rect 13354 5148 13360 5160
rect 13315 5120 13360 5148
rect 13354 5108 13360 5120
rect 13412 5108 13418 5160
rect 17402 5108 17408 5160
rect 17460 5148 17466 5160
rect 17569 5151 17627 5157
rect 17569 5148 17581 5151
rect 17460 5120 17581 5148
rect 17460 5108 17466 5120
rect 17569 5117 17581 5120
rect 17615 5117 17627 5151
rect 17569 5111 17627 5117
rect 20625 5151 20683 5157
rect 20625 5117 20637 5151
rect 20671 5117 20683 5151
rect 21358 5148 21364 5160
rect 21319 5120 21364 5148
rect 20625 5111 20683 5117
rect 9272 5052 9628 5080
rect 15841 5083 15899 5089
rect 9272 5040 9278 5052
rect 15841 5049 15853 5083
rect 15887 5080 15899 5083
rect 16482 5080 16488 5092
rect 15887 5052 16488 5080
rect 15887 5049 15899 5052
rect 15841 5043 15899 5049
rect 16482 5040 16488 5052
rect 16540 5040 16546 5092
rect 20640 5080 20668 5111
rect 21358 5108 21364 5120
rect 21416 5108 21422 5160
rect 22741 5151 22799 5157
rect 22741 5117 22753 5151
rect 22787 5117 22799 5151
rect 22741 5111 22799 5117
rect 21453 5083 21511 5089
rect 21453 5080 21465 5083
rect 20640 5052 21465 5080
rect 21453 5049 21465 5052
rect 21499 5049 21511 5083
rect 22756 5080 22784 5111
rect 22922 5108 22928 5160
rect 22980 5148 22986 5160
rect 23216 5157 23244 5188
rect 23201 5151 23259 5157
rect 23201 5148 23213 5151
rect 22980 5120 23213 5148
rect 22980 5108 22986 5120
rect 23201 5117 23213 5120
rect 23247 5117 23259 5151
rect 23201 5111 23259 5117
rect 23385 5151 23443 5157
rect 23385 5117 23397 5151
rect 23431 5148 23443 5151
rect 23474 5148 23480 5160
rect 23431 5120 23480 5148
rect 23431 5117 23443 5120
rect 23385 5111 23443 5117
rect 23400 5080 23428 5111
rect 23474 5108 23480 5120
rect 23532 5108 23538 5160
rect 24136 5157 24164 5188
rect 25958 5176 25964 5188
rect 26016 5176 26022 5228
rect 26068 5225 26096 5256
rect 30929 5253 30941 5287
rect 30975 5284 30987 5287
rect 31294 5284 31300 5296
rect 30975 5256 31300 5284
rect 30975 5253 30987 5256
rect 30929 5247 30987 5253
rect 31294 5244 31300 5256
rect 31352 5244 31358 5296
rect 26053 5219 26111 5225
rect 26053 5185 26065 5219
rect 26099 5185 26111 5219
rect 32306 5216 32312 5228
rect 26053 5179 26111 5185
rect 31220 5188 32312 5216
rect 24121 5151 24179 5157
rect 24121 5117 24133 5151
rect 24167 5117 24179 5151
rect 24121 5111 24179 5117
rect 24302 5108 24308 5160
rect 24360 5148 24366 5160
rect 25976 5148 26004 5176
rect 24360 5120 26004 5148
rect 30193 5151 30251 5157
rect 24360 5108 24366 5120
rect 30193 5117 30205 5151
rect 30239 5117 30251 5151
rect 30374 5148 30380 5160
rect 30335 5120 30380 5148
rect 30193 5111 30251 5117
rect 22756 5052 23428 5080
rect 30208 5080 30236 5111
rect 30374 5108 30380 5120
rect 30432 5108 30438 5160
rect 31220 5157 31248 5188
rect 32306 5176 32312 5188
rect 32364 5176 32370 5228
rect 31021 5151 31079 5157
rect 31021 5117 31033 5151
rect 31067 5117 31079 5151
rect 31021 5111 31079 5117
rect 31205 5151 31263 5157
rect 31205 5117 31217 5151
rect 31251 5117 31263 5151
rect 31662 5148 31668 5160
rect 31623 5120 31668 5148
rect 31205 5111 31263 5117
rect 31036 5080 31064 5111
rect 31662 5108 31668 5120
rect 31720 5108 31726 5160
rect 31938 5148 31944 5160
rect 31851 5120 31944 5148
rect 31938 5108 31944 5120
rect 31996 5148 32002 5160
rect 32950 5148 32956 5160
rect 31996 5120 32956 5148
rect 31996 5108 32002 5120
rect 32950 5108 32956 5120
rect 33008 5108 33014 5160
rect 33042 5108 33048 5160
rect 33100 5148 33106 5160
rect 33413 5151 33471 5157
rect 33413 5148 33425 5151
rect 33100 5120 33425 5148
rect 33100 5108 33106 5120
rect 33413 5117 33425 5120
rect 33459 5117 33471 5151
rect 33413 5111 33471 5117
rect 31478 5080 31484 5092
rect 30208 5052 31484 5080
rect 21453 5043 21511 5049
rect 31478 5040 31484 5052
rect 31536 5040 31542 5092
rect 5534 4972 5540 5024
rect 5592 5012 5598 5024
rect 5592 4984 5637 5012
rect 5592 4972 5598 4984
rect 15010 4972 15016 5024
rect 15068 5012 15074 5024
rect 15473 5015 15531 5021
rect 15473 5012 15485 5015
rect 15068 4984 15485 5012
rect 15068 4972 15074 4984
rect 15473 4981 15485 4984
rect 15519 4981 15531 5015
rect 15473 4975 15531 4981
rect 15933 5015 15991 5021
rect 15933 4981 15945 5015
rect 15979 5012 15991 5015
rect 16114 5012 16120 5024
rect 15979 4984 16120 5012
rect 15979 4981 15991 4984
rect 15933 4975 15991 4981
rect 16114 4972 16120 4984
rect 16172 4972 16178 5024
rect 17954 4972 17960 5024
rect 18012 5012 18018 5024
rect 18693 5015 18751 5021
rect 18693 5012 18705 5015
rect 18012 4984 18705 5012
rect 18012 4972 18018 4984
rect 18693 4981 18705 4984
rect 18739 4981 18751 5015
rect 20898 5012 20904 5024
rect 20859 4984 20904 5012
rect 18693 4975 18751 4981
rect 20898 4972 20904 4984
rect 20956 4972 20962 5024
rect 25869 5015 25927 5021
rect 25869 4981 25881 5015
rect 25915 5012 25927 5015
rect 27062 5012 27068 5024
rect 25915 4984 27068 5012
rect 25915 4981 25927 4984
rect 25869 4975 25927 4981
rect 27062 4972 27068 4984
rect 27120 4972 27126 5024
rect 30285 5015 30343 5021
rect 30285 4981 30297 5015
rect 30331 5012 30343 5015
rect 30558 5012 30564 5024
rect 30331 4984 30564 5012
rect 30331 4981 30343 4984
rect 30285 4975 30343 4981
rect 30558 4972 30564 4984
rect 30616 4972 30622 5024
rect 31757 5015 31815 5021
rect 31757 4981 31769 5015
rect 31803 5012 31815 5015
rect 31846 5012 31852 5024
rect 31803 4984 31852 5012
rect 31803 4981 31815 4984
rect 31757 4975 31815 4981
rect 31846 4972 31852 4984
rect 31904 4972 31910 5024
rect 33410 4972 33416 5024
rect 33468 5012 33474 5024
rect 33505 5015 33563 5021
rect 33505 5012 33517 5015
rect 33468 4984 33517 5012
rect 33468 4972 33474 4984
rect 33505 4981 33517 4984
rect 33551 4981 33563 5015
rect 33505 4975 33563 4981
rect 1104 4922 34316 4944
rect 1104 4870 12052 4922
rect 12104 4870 12116 4922
rect 12168 4870 12180 4922
rect 12232 4870 12244 4922
rect 12296 4870 23123 4922
rect 23175 4870 23187 4922
rect 23239 4870 23251 4922
rect 23303 4870 23315 4922
rect 23367 4870 34316 4922
rect 1104 4848 34316 4870
rect 12986 4808 12992 4820
rect 2746 4780 12992 4808
rect 1949 4743 2007 4749
rect 1949 4709 1961 4743
rect 1995 4740 2007 4743
rect 2746 4740 2774 4780
rect 12986 4768 12992 4780
rect 13044 4768 13050 4820
rect 13722 4768 13728 4820
rect 13780 4808 13786 4820
rect 13780 4780 15516 4808
rect 13780 4768 13786 4780
rect 1995 4712 2774 4740
rect 2961 4743 3019 4749
rect 1995 4709 2007 4712
rect 1949 4703 2007 4709
rect 2961 4709 2973 4743
rect 3007 4740 3019 4743
rect 3050 4740 3056 4752
rect 3007 4712 3056 4740
rect 3007 4709 3019 4712
rect 2961 4703 3019 4709
rect 3050 4700 3056 4712
rect 3108 4700 3114 4752
rect 5166 4700 5172 4752
rect 5224 4700 5230 4752
rect 15010 4740 15016 4752
rect 14971 4712 15016 4740
rect 15010 4700 15016 4712
rect 15068 4700 15074 4752
rect 15488 4726 15516 4780
rect 17310 4768 17316 4820
rect 17368 4808 17374 4820
rect 17773 4811 17831 4817
rect 17773 4808 17785 4811
rect 17368 4780 17785 4808
rect 17368 4768 17374 4780
rect 17773 4777 17785 4780
rect 17819 4777 17831 4811
rect 22370 4808 22376 4820
rect 22283 4780 22376 4808
rect 17773 4771 17831 4777
rect 22370 4768 22376 4780
rect 22428 4808 22434 4820
rect 23293 4811 23351 4817
rect 23293 4808 23305 4811
rect 22428 4780 23305 4808
rect 22428 4768 22434 4780
rect 23293 4777 23305 4780
rect 23339 4777 23351 4811
rect 23293 4771 23351 4777
rect 31846 4768 31852 4820
rect 31904 4808 31910 4820
rect 31941 4811 31999 4817
rect 31941 4808 31953 4811
rect 31904 4780 31953 4808
rect 31904 4768 31910 4780
rect 31941 4777 31953 4780
rect 31987 4777 31999 4811
rect 31941 4771 31999 4777
rect 16298 4700 16304 4752
rect 16356 4740 16362 4752
rect 16356 4712 20300 4740
rect 16356 4700 16362 4712
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 4522 4672 4528 4684
rect 4295 4644 4528 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 4522 4632 4528 4644
rect 4580 4632 4586 4684
rect 14734 4672 14740 4684
rect 14695 4644 14740 4672
rect 14734 4632 14740 4644
rect 14792 4632 14798 4684
rect 17773 4675 17831 4681
rect 17773 4641 17785 4675
rect 17819 4641 17831 4675
rect 17954 4672 17960 4684
rect 17915 4644 17960 4672
rect 17773 4635 17831 4641
rect 3050 4604 3056 4616
rect 3011 4576 3056 4604
rect 3050 4564 3056 4576
rect 3108 4564 3114 4616
rect 3234 4604 3240 4616
rect 3195 4576 3240 4604
rect 3234 4564 3240 4576
rect 3292 4564 3298 4616
rect 4614 4604 4620 4616
rect 4575 4576 4620 4604
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 17788 4536 17816 4635
rect 17954 4632 17960 4644
rect 18012 4632 18018 4684
rect 18322 4632 18328 4684
rect 18380 4672 18386 4684
rect 18785 4675 18843 4681
rect 18785 4672 18797 4675
rect 18380 4644 18797 4672
rect 18380 4632 18386 4644
rect 18785 4641 18797 4644
rect 18831 4641 18843 4675
rect 18785 4635 18843 4641
rect 18877 4675 18935 4681
rect 18877 4641 18889 4675
rect 18923 4672 18935 4675
rect 19150 4672 19156 4684
rect 18923 4644 19156 4672
rect 18923 4641 18935 4644
rect 18877 4635 18935 4641
rect 19150 4632 19156 4644
rect 19208 4632 19214 4684
rect 19886 4632 19892 4684
rect 19944 4672 19950 4684
rect 19981 4675 20039 4681
rect 19981 4672 19993 4675
rect 19944 4644 19993 4672
rect 19944 4632 19950 4644
rect 19981 4641 19993 4644
rect 20027 4641 20039 4675
rect 20162 4672 20168 4684
rect 20123 4644 20168 4672
rect 19981 4635 20039 4641
rect 20162 4632 20168 4644
rect 20220 4632 20226 4684
rect 20272 4672 20300 4712
rect 20898 4700 20904 4752
rect 20956 4740 20962 4752
rect 21238 4743 21296 4749
rect 21238 4740 21250 4743
rect 20956 4712 21250 4740
rect 20956 4700 20962 4712
rect 21238 4709 21250 4712
rect 21284 4709 21296 4743
rect 28074 4740 28080 4752
rect 21238 4703 21296 4709
rect 27448 4712 28080 4740
rect 23201 4675 23259 4681
rect 20272 4644 22094 4672
rect 19061 4607 19119 4613
rect 19061 4573 19073 4607
rect 19107 4604 19119 4607
rect 20073 4607 20131 4613
rect 20073 4604 20085 4607
rect 19107 4576 20085 4604
rect 19107 4573 19119 4576
rect 19061 4567 19119 4573
rect 20073 4573 20085 4576
rect 20119 4573 20131 4607
rect 20073 4567 20131 4573
rect 20714 4564 20720 4616
rect 20772 4604 20778 4616
rect 20993 4607 21051 4613
rect 20993 4604 21005 4607
rect 20772 4576 21005 4604
rect 20772 4564 20778 4576
rect 20993 4573 21005 4576
rect 21039 4573 21051 4607
rect 22066 4604 22094 4644
rect 23201 4641 23213 4675
rect 23247 4672 23259 4675
rect 24394 4672 24400 4684
rect 23247 4644 24400 4672
rect 23247 4641 23259 4644
rect 23201 4635 23259 4641
rect 24394 4632 24400 4644
rect 24452 4632 24458 4684
rect 27448 4681 27476 4712
rect 28074 4700 28080 4712
rect 28132 4740 28138 4752
rect 28534 4740 28540 4752
rect 28132 4712 28540 4740
rect 28132 4700 28138 4712
rect 28534 4700 28540 4712
rect 28592 4700 28598 4752
rect 30653 4743 30711 4749
rect 30653 4709 30665 4743
rect 30699 4740 30711 4743
rect 31297 4743 31355 4749
rect 31297 4740 31309 4743
rect 30699 4712 31309 4740
rect 30699 4709 30711 4712
rect 30653 4703 30711 4709
rect 31297 4709 31309 4712
rect 31343 4740 31355 4743
rect 33410 4740 33416 4752
rect 31343 4712 31984 4740
rect 33371 4712 33416 4740
rect 31343 4709 31355 4712
rect 31297 4703 31355 4709
rect 27433 4675 27491 4681
rect 27433 4641 27445 4675
rect 27479 4641 27491 4675
rect 27614 4672 27620 4684
rect 27575 4644 27620 4672
rect 27433 4635 27491 4641
rect 27614 4632 27620 4644
rect 27672 4632 27678 4684
rect 27709 4675 27767 4681
rect 27709 4641 27721 4675
rect 27755 4672 27767 4675
rect 28442 4672 28448 4684
rect 27755 4644 28448 4672
rect 27755 4641 27767 4644
rect 27709 4635 27767 4641
rect 28442 4632 28448 4644
rect 28500 4632 28506 4684
rect 30558 4672 30564 4684
rect 30519 4644 30564 4672
rect 30558 4632 30564 4644
rect 30616 4632 30622 4684
rect 30742 4672 30748 4684
rect 30703 4644 30748 4672
rect 30742 4632 30748 4644
rect 30800 4632 30806 4684
rect 31202 4672 31208 4684
rect 31163 4644 31208 4672
rect 31202 4632 31208 4644
rect 31260 4632 31266 4684
rect 31481 4675 31539 4681
rect 31481 4641 31493 4675
rect 31527 4672 31539 4675
rect 31846 4672 31852 4684
rect 31527 4644 31852 4672
rect 31527 4641 31539 4644
rect 31481 4635 31539 4641
rect 31846 4632 31852 4644
rect 31904 4632 31910 4684
rect 31956 4681 31984 4712
rect 33410 4700 33416 4712
rect 33468 4700 33474 4752
rect 33594 4740 33600 4752
rect 33555 4712 33600 4740
rect 33594 4700 33600 4712
rect 33652 4700 33658 4752
rect 31941 4675 31999 4681
rect 31941 4641 31953 4675
rect 31987 4641 31999 4675
rect 31941 4635 31999 4641
rect 32125 4675 32183 4681
rect 32125 4641 32137 4675
rect 32171 4672 32183 4675
rect 32306 4672 32312 4684
rect 32171 4644 32312 4672
rect 32171 4641 32183 4644
rect 32125 4635 32183 4641
rect 32306 4632 32312 4644
rect 32364 4632 32370 4684
rect 23385 4607 23443 4613
rect 23385 4604 23397 4607
rect 22066 4576 23397 4604
rect 20993 4567 21051 4573
rect 23385 4573 23397 4576
rect 23431 4604 23443 4607
rect 25682 4604 25688 4616
rect 23431 4576 25688 4604
rect 23431 4573 23443 4576
rect 23385 4567 23443 4573
rect 25682 4564 25688 4576
rect 25740 4564 25746 4616
rect 29454 4564 29460 4616
rect 29512 4604 29518 4616
rect 33042 4604 33048 4616
rect 29512 4576 33048 4604
rect 29512 4564 29518 4576
rect 33042 4564 33048 4576
rect 33100 4564 33106 4616
rect 20622 4536 20628 4548
rect 17788 4508 20628 4536
rect 20622 4496 20628 4508
rect 20680 4536 20686 4548
rect 20680 4508 21036 4536
rect 20680 4496 20686 4508
rect 21008 4480 21036 4508
rect 27062 4496 27068 4548
rect 27120 4536 27126 4548
rect 32490 4536 32496 4548
rect 27120 4508 32496 4536
rect 27120 4496 27126 4508
rect 32490 4496 32496 4508
rect 32548 4496 32554 4548
rect 1854 4468 1860 4480
rect 1815 4440 1860 4468
rect 1854 4428 1860 4440
rect 1912 4428 1918 4480
rect 2590 4468 2596 4480
rect 2551 4440 2596 4468
rect 2590 4428 2596 4440
rect 2648 4428 2654 4480
rect 5626 4428 5632 4480
rect 5684 4468 5690 4480
rect 6043 4471 6101 4477
rect 6043 4468 6055 4471
rect 5684 4440 6055 4468
rect 5684 4428 5690 4440
rect 6043 4437 6055 4440
rect 6089 4437 6101 4471
rect 16482 4468 16488 4480
rect 16443 4440 16488 4468
rect 6043 4431 6101 4437
rect 16482 4428 16488 4440
rect 16540 4428 16546 4480
rect 18966 4428 18972 4480
rect 19024 4468 19030 4480
rect 19024 4440 19069 4468
rect 19024 4428 19030 4440
rect 20990 4428 20996 4480
rect 21048 4428 21054 4480
rect 22833 4471 22891 4477
rect 22833 4437 22845 4471
rect 22879 4468 22891 4471
rect 22922 4468 22928 4480
rect 22879 4440 22928 4468
rect 22879 4437 22891 4440
rect 22833 4431 22891 4437
rect 22922 4428 22928 4440
rect 22980 4428 22986 4480
rect 26786 4428 26792 4480
rect 26844 4468 26850 4480
rect 27249 4471 27307 4477
rect 27249 4468 27261 4471
rect 26844 4440 27261 4468
rect 26844 4428 26850 4440
rect 27249 4437 27261 4440
rect 27295 4437 27307 4471
rect 27249 4431 27307 4437
rect 31481 4471 31539 4477
rect 31481 4437 31493 4471
rect 31527 4468 31539 4471
rect 31846 4468 31852 4480
rect 31527 4440 31852 4468
rect 31527 4437 31539 4440
rect 31481 4431 31539 4437
rect 31846 4428 31852 4440
rect 31904 4428 31910 4480
rect 1104 4378 34316 4400
rect 1104 4326 6517 4378
rect 6569 4326 6581 4378
rect 6633 4326 6645 4378
rect 6697 4326 6709 4378
rect 6761 4326 17588 4378
rect 17640 4326 17652 4378
rect 17704 4326 17716 4378
rect 17768 4326 17780 4378
rect 17832 4326 28658 4378
rect 28710 4326 28722 4378
rect 28774 4326 28786 4378
rect 28838 4326 28850 4378
rect 28902 4326 34316 4378
rect 1104 4304 34316 4326
rect 3050 4224 3056 4276
rect 3108 4264 3114 4276
rect 3743 4267 3801 4273
rect 3743 4264 3755 4267
rect 3108 4236 3755 4264
rect 3108 4224 3114 4236
rect 3743 4233 3755 4236
rect 3789 4264 3801 4267
rect 4062 4264 4068 4276
rect 3789 4236 4068 4264
rect 3789 4233 3801 4236
rect 3743 4227 3801 4233
rect 4062 4224 4068 4236
rect 4120 4224 4126 4276
rect 9582 4273 9588 4276
rect 9572 4267 9588 4273
rect 9572 4233 9584 4267
rect 9572 4227 9588 4233
rect 9582 4224 9588 4227
rect 9640 4224 9646 4276
rect 14479 4267 14537 4273
rect 14479 4233 14491 4267
rect 14525 4264 14537 4267
rect 14642 4264 14648 4276
rect 14525 4236 14648 4264
rect 14525 4233 14537 4236
rect 14479 4227 14537 4233
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 20806 4224 20812 4276
rect 20864 4264 20870 4276
rect 22922 4273 22928 4276
rect 20901 4267 20959 4273
rect 20901 4264 20913 4267
rect 20864 4236 20913 4264
rect 20864 4224 20870 4236
rect 20901 4233 20913 4236
rect 20947 4233 20959 4267
rect 20901 4227 20959 4233
rect 22912 4267 22928 4273
rect 22912 4233 22924 4267
rect 22912 4227 22928 4233
rect 22922 4224 22928 4227
rect 22980 4224 22986 4276
rect 27614 4224 27620 4276
rect 27672 4264 27678 4276
rect 28077 4267 28135 4273
rect 28077 4264 28089 4267
rect 27672 4236 28089 4264
rect 27672 4224 27678 4236
rect 28077 4233 28089 4236
rect 28123 4233 28135 4267
rect 28077 4227 28135 4233
rect 28442 4224 28448 4276
rect 28500 4264 28506 4276
rect 29454 4264 29460 4276
rect 28500 4236 29460 4264
rect 28500 4224 28506 4236
rect 29454 4224 29460 4236
rect 29512 4224 29518 4276
rect 31202 4224 31208 4276
rect 31260 4264 31266 4276
rect 31389 4267 31447 4273
rect 31389 4264 31401 4267
rect 31260 4236 31401 4264
rect 31260 4224 31266 4236
rect 31389 4233 31401 4236
rect 31435 4233 31447 4267
rect 31389 4227 31447 4233
rect 29086 4196 29092 4208
rect 28460 4168 29092 4196
rect 1394 4088 1400 4140
rect 1452 4128 1458 4140
rect 1949 4131 2007 4137
rect 1949 4128 1961 4131
rect 1452 4100 1961 4128
rect 1452 4088 1458 4100
rect 1949 4097 1961 4100
rect 1995 4097 2007 4131
rect 1949 4091 2007 4097
rect 2317 4131 2375 4137
rect 2317 4097 2329 4131
rect 2363 4128 2375 4131
rect 2590 4128 2596 4140
rect 2363 4100 2596 4128
rect 2363 4097 2375 4100
rect 2317 4091 2375 4097
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 5350 4128 5356 4140
rect 5311 4100 5356 4128
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 5445 4131 5503 4137
rect 5445 4097 5457 4131
rect 5491 4128 5503 4131
rect 5534 4128 5540 4140
rect 5491 4100 5540 4128
rect 5491 4097 5503 4100
rect 5445 4091 5503 4097
rect 5534 4088 5540 4100
rect 5592 4088 5598 4140
rect 9306 4128 9312 4140
rect 9267 4100 9312 4128
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 10318 4088 10324 4140
rect 10376 4128 10382 4140
rect 11057 4131 11115 4137
rect 11057 4128 11069 4131
rect 10376 4100 11069 4128
rect 10376 4088 10382 4100
rect 11057 4097 11069 4100
rect 11103 4097 11115 4131
rect 12986 4128 12992 4140
rect 12947 4100 12992 4128
rect 11057 4091 11115 4097
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 14734 4128 14740 4140
rect 14695 4100 14740 4128
rect 14734 4088 14740 4100
rect 14792 4088 14798 4140
rect 17126 4088 17132 4140
rect 17184 4128 17190 4140
rect 18877 4131 18935 4137
rect 18877 4128 18889 4131
rect 17184 4100 18889 4128
rect 17184 4088 17190 4100
rect 18877 4097 18889 4100
rect 18923 4097 18935 4131
rect 21082 4128 21088 4140
rect 18877 4091 18935 4097
rect 20824 4100 21088 4128
rect 18966 4020 18972 4072
rect 19024 4060 19030 4072
rect 20824 4069 20852 4100
rect 21082 4088 21088 4100
rect 21140 4128 21146 4140
rect 22370 4128 22376 4140
rect 21140 4100 22376 4128
rect 21140 4088 21146 4100
rect 22370 4088 22376 4100
rect 22428 4088 22434 4140
rect 28460 4137 28488 4168
rect 29086 4156 29092 4168
rect 29144 4156 29150 4208
rect 29196 4168 30512 4196
rect 28445 4131 28503 4137
rect 28445 4097 28457 4131
rect 28491 4097 28503 4131
rect 29196 4128 29224 4168
rect 28445 4091 28503 4097
rect 28552 4100 29224 4128
rect 28552 4072 28580 4100
rect 19133 4063 19191 4069
rect 19133 4060 19145 4063
rect 19024 4032 19145 4060
rect 19024 4020 19030 4032
rect 19133 4029 19145 4032
rect 19179 4029 19191 4063
rect 19133 4023 19191 4029
rect 20809 4063 20867 4069
rect 20809 4029 20821 4063
rect 20855 4029 20867 4063
rect 20990 4060 20996 4072
rect 20951 4032 20996 4060
rect 20809 4023 20867 4029
rect 20990 4020 20996 4032
rect 21048 4020 21054 4072
rect 22649 4063 22707 4069
rect 22649 4060 22661 4063
rect 22066 4032 22661 4060
rect 5166 3992 5172 4004
rect 3358 3964 5172 3992
rect 5166 3952 5172 3964
rect 5224 3952 5230 4004
rect 5537 3995 5595 4001
rect 5537 3961 5549 3995
rect 5583 3992 5595 3995
rect 5626 3992 5632 4004
rect 5583 3964 5632 3992
rect 5583 3961 5595 3964
rect 5537 3955 5595 3961
rect 5626 3952 5632 3964
rect 5684 3952 5690 4004
rect 10810 3964 12434 3992
rect 5905 3927 5963 3933
rect 5905 3893 5917 3927
rect 5951 3924 5963 3927
rect 7006 3924 7012 3936
rect 5951 3896 7012 3924
rect 5951 3893 5963 3896
rect 5905 3887 5963 3893
rect 7006 3884 7012 3896
rect 7064 3884 7070 3936
rect 12406 3924 12434 3964
rect 13722 3952 13728 4004
rect 13780 3952 13786 4004
rect 20714 3952 20720 4004
rect 20772 3992 20778 4004
rect 22066 3992 22094 4032
rect 22649 4029 22661 4032
rect 22695 4029 22707 4063
rect 27522 4060 27528 4072
rect 24058 4032 27528 4060
rect 22649 4023 22707 4029
rect 27522 4020 27528 4032
rect 27580 4020 27586 4072
rect 28353 4063 28411 4069
rect 28353 4029 28365 4063
rect 28399 4060 28411 4063
rect 28534 4060 28540 4072
rect 28399 4032 28540 4060
rect 28399 4029 28411 4032
rect 28353 4023 28411 4029
rect 28534 4020 28540 4032
rect 28592 4020 28598 4072
rect 28626 4020 28632 4072
rect 28684 4060 28690 4072
rect 29181 4063 29239 4069
rect 29181 4060 29193 4063
rect 28684 4032 29193 4060
rect 28684 4020 28690 4032
rect 29181 4029 29193 4032
rect 29227 4029 29239 4063
rect 29454 4060 29460 4072
rect 29415 4032 29460 4060
rect 29181 4023 29239 4029
rect 29454 4020 29460 4032
rect 29512 4020 29518 4072
rect 30282 4060 30288 4072
rect 30243 4032 30288 4060
rect 30282 4020 30288 4032
rect 30340 4020 30346 4072
rect 30484 4069 30512 4168
rect 30742 4156 30748 4208
rect 30800 4156 30806 4208
rect 30653 4131 30711 4137
rect 30653 4097 30665 4131
rect 30699 4128 30711 4131
rect 30760 4128 30788 4156
rect 31478 4128 31484 4140
rect 30699 4100 30788 4128
rect 31439 4100 31484 4128
rect 30699 4097 30711 4100
rect 30653 4091 30711 4097
rect 31478 4088 31484 4100
rect 31536 4088 31542 4140
rect 30469 4063 30527 4069
rect 30469 4029 30481 4063
rect 30515 4060 30527 4063
rect 30742 4060 30748 4072
rect 30515 4032 30748 4060
rect 30515 4029 30527 4032
rect 30469 4023 30527 4029
rect 30742 4020 30748 4032
rect 30800 4020 30806 4072
rect 31202 4060 31208 4072
rect 31163 4032 31208 4060
rect 31202 4020 31208 4032
rect 31260 4020 31266 4072
rect 31297 4063 31355 4069
rect 31297 4029 31309 4063
rect 31343 4029 31355 4063
rect 31297 4023 31355 4029
rect 28442 3992 28448 4004
rect 20772 3964 22094 3992
rect 24320 3964 28448 3992
rect 20772 3952 20778 3964
rect 13740 3924 13768 3952
rect 12406 3896 13768 3924
rect 20162 3884 20168 3936
rect 20220 3924 20226 3936
rect 20257 3927 20315 3933
rect 20257 3924 20269 3927
rect 20220 3896 20269 3924
rect 20220 3884 20226 3896
rect 20257 3893 20269 3896
rect 20303 3924 20315 3927
rect 24320 3924 24348 3964
rect 28442 3952 28448 3964
rect 28500 3952 28506 4004
rect 30374 3992 30380 4004
rect 28552 3964 30380 3992
rect 20303 3896 24348 3924
rect 20303 3893 20315 3896
rect 20257 3887 20315 3893
rect 24394 3884 24400 3936
rect 24452 3924 24458 3936
rect 28552 3924 28580 3964
rect 30374 3952 30380 3964
rect 30432 3952 30438 4004
rect 31312 3992 31340 4023
rect 31220 3964 31340 3992
rect 24452 3896 28580 3924
rect 28997 3927 29055 3933
rect 24452 3884 24458 3896
rect 28997 3893 29009 3927
rect 29043 3924 29055 3927
rect 29086 3924 29092 3936
rect 29043 3896 29092 3924
rect 29043 3893 29055 3896
rect 28997 3887 29055 3893
rect 29086 3884 29092 3896
rect 29144 3884 29150 3936
rect 29365 3927 29423 3933
rect 29365 3893 29377 3927
rect 29411 3924 29423 3927
rect 29546 3924 29552 3936
rect 29411 3896 29552 3924
rect 29411 3893 29423 3896
rect 29365 3887 29423 3893
rect 29546 3884 29552 3896
rect 29604 3884 29610 3936
rect 30190 3884 30196 3936
rect 30248 3924 30254 3936
rect 31220 3924 31248 3964
rect 30248 3896 31248 3924
rect 30248 3884 30254 3896
rect 1104 3834 34316 3856
rect 1104 3782 12052 3834
rect 12104 3782 12116 3834
rect 12168 3782 12180 3834
rect 12232 3782 12244 3834
rect 12296 3782 23123 3834
rect 23175 3782 23187 3834
rect 23239 3782 23251 3834
rect 23303 3782 23315 3834
rect 23367 3782 34316 3834
rect 1104 3760 34316 3782
rect 4249 3723 4307 3729
rect 4249 3689 4261 3723
rect 4295 3720 4307 3723
rect 4614 3720 4620 3732
rect 4295 3692 4620 3720
rect 4295 3689 4307 3692
rect 4249 3683 4307 3689
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 5534 3680 5540 3732
rect 5592 3729 5598 3732
rect 5592 3723 5641 3729
rect 5592 3689 5595 3723
rect 5629 3689 5641 3723
rect 5592 3683 5641 3689
rect 5592 3680 5598 3683
rect 6914 3680 6920 3732
rect 6972 3720 6978 3732
rect 29546 3720 29552 3732
rect 6972 3692 7420 3720
rect 29507 3692 29552 3720
rect 6972 3680 6978 3692
rect 5166 3612 5172 3664
rect 5224 3652 5230 3664
rect 5224 3624 6026 3652
rect 5224 3612 5230 3624
rect 4062 3544 4068 3596
rect 4120 3584 4126 3596
rect 4617 3587 4675 3593
rect 4617 3584 4629 3587
rect 4120 3556 4629 3584
rect 4120 3544 4126 3556
rect 4617 3553 4629 3556
rect 4663 3553 4675 3587
rect 4617 3547 4675 3553
rect 4709 3587 4767 3593
rect 4709 3553 4721 3587
rect 4755 3584 4767 3587
rect 5626 3584 5632 3596
rect 4755 3556 5632 3584
rect 4755 3553 4767 3556
rect 4709 3547 4767 3553
rect 5626 3544 5632 3556
rect 5684 3544 5690 3596
rect 7006 3584 7012 3596
rect 6967 3556 7012 3584
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 7392 3593 7420 3692
rect 29546 3680 29552 3692
rect 29604 3680 29610 3732
rect 31478 3680 31484 3732
rect 31536 3720 31542 3732
rect 33321 3723 33379 3729
rect 33321 3720 33333 3723
rect 31536 3692 33333 3720
rect 31536 3680 31542 3692
rect 33321 3689 33333 3692
rect 33367 3689 33379 3723
rect 33321 3683 33379 3689
rect 17126 3612 17132 3664
rect 17184 3652 17190 3664
rect 26786 3652 26792 3664
rect 17184 3624 17540 3652
rect 26747 3624 26792 3652
rect 17184 3612 17190 3624
rect 7377 3587 7435 3593
rect 7377 3553 7389 3587
rect 7423 3553 7435 3587
rect 7377 3547 7435 3553
rect 17241 3587 17299 3593
rect 17241 3553 17253 3587
rect 17287 3584 17299 3587
rect 17402 3584 17408 3596
rect 17287 3556 17408 3584
rect 17287 3553 17299 3556
rect 17241 3547 17299 3553
rect 17402 3544 17408 3556
rect 17460 3544 17466 3596
rect 17512 3593 17540 3624
rect 26786 3612 26792 3624
rect 26844 3612 26850 3664
rect 27522 3612 27528 3664
rect 27580 3612 27586 3664
rect 28534 3652 28540 3664
rect 28495 3624 28540 3652
rect 28534 3612 28540 3624
rect 28592 3612 28598 3664
rect 31202 3652 31208 3664
rect 29380 3624 31208 3652
rect 17497 3587 17555 3593
rect 17497 3553 17509 3587
rect 17543 3553 17555 3587
rect 18138 3584 18144 3596
rect 18099 3556 18144 3584
rect 17497 3547 17555 3553
rect 18138 3544 18144 3556
rect 18196 3544 18202 3596
rect 18233 3587 18291 3593
rect 18233 3553 18245 3587
rect 18279 3584 18291 3587
rect 19150 3584 19156 3596
rect 18279 3556 19156 3584
rect 18279 3553 18291 3556
rect 18233 3547 18291 3553
rect 19150 3544 19156 3556
rect 19208 3544 19214 3596
rect 20993 3587 21051 3593
rect 20993 3553 21005 3587
rect 21039 3584 21051 3587
rect 21082 3584 21088 3596
rect 21039 3556 21088 3584
rect 21039 3553 21051 3556
rect 20993 3547 21051 3553
rect 21082 3544 21088 3556
rect 21140 3544 21146 3596
rect 29178 3544 29184 3596
rect 29236 3584 29242 3596
rect 29380 3593 29408 3624
rect 31202 3612 31208 3624
rect 31260 3612 31266 3664
rect 31846 3652 31852 3664
rect 31807 3624 31852 3652
rect 31846 3612 31852 3624
rect 31904 3612 31910 3664
rect 32858 3612 32864 3664
rect 32916 3612 32922 3664
rect 29273 3587 29331 3593
rect 29273 3584 29285 3587
rect 29236 3556 29285 3584
rect 29236 3544 29242 3556
rect 29273 3553 29285 3556
rect 29319 3553 29331 3587
rect 29273 3547 29331 3553
rect 29365 3587 29423 3593
rect 29365 3553 29377 3587
rect 29411 3553 29423 3587
rect 30742 3584 30748 3596
rect 30703 3556 30748 3584
rect 29365 3547 29423 3553
rect 4893 3519 4951 3525
rect 4893 3485 4905 3519
rect 4939 3516 4951 3519
rect 5350 3516 5356 3528
rect 4939 3488 5356 3516
rect 4939 3485 4951 3488
rect 4893 3479 4951 3485
rect 5350 3476 5356 3488
rect 5408 3476 5414 3528
rect 18414 3516 18420 3528
rect 18375 3488 18420 3516
rect 18414 3476 18420 3488
rect 18472 3476 18478 3528
rect 26510 3516 26516 3528
rect 26471 3488 26516 3516
rect 26510 3476 26516 3488
rect 26568 3476 26574 3528
rect 16114 3380 16120 3392
rect 16075 3352 16120 3380
rect 16114 3340 16120 3352
rect 16172 3340 16178 3392
rect 18322 3340 18328 3392
rect 18380 3380 18386 3392
rect 18380 3352 18425 3380
rect 18380 3340 18386 3352
rect 20438 3340 20444 3392
rect 20496 3380 20502 3392
rect 20901 3383 20959 3389
rect 20901 3380 20913 3383
rect 20496 3352 20913 3380
rect 20496 3340 20502 3352
rect 20901 3349 20913 3352
rect 20947 3349 20959 3383
rect 29288 3380 29316 3547
rect 30742 3544 30748 3556
rect 30800 3544 30806 3596
rect 31570 3584 31576 3596
rect 31531 3556 31576 3584
rect 31570 3544 31576 3556
rect 31628 3544 31634 3596
rect 29549 3519 29607 3525
rect 29549 3485 29561 3519
rect 29595 3485 29607 3519
rect 29549 3479 29607 3485
rect 29564 3448 29592 3479
rect 30282 3476 30288 3528
rect 30340 3516 30346 3528
rect 30469 3519 30527 3525
rect 30469 3516 30481 3519
rect 30340 3488 30481 3516
rect 30340 3476 30346 3488
rect 30469 3485 30481 3488
rect 30515 3485 30527 3519
rect 30469 3479 30527 3485
rect 30561 3451 30619 3457
rect 30561 3448 30573 3451
rect 29564 3420 30573 3448
rect 30561 3417 30573 3420
rect 30607 3417 30619 3451
rect 30561 3411 30619 3417
rect 30190 3380 30196 3392
rect 29288 3352 30196 3380
rect 20901 3343 20959 3349
rect 30190 3340 30196 3352
rect 30248 3380 30254 3392
rect 30653 3383 30711 3389
rect 30653 3380 30665 3383
rect 30248 3352 30665 3380
rect 30248 3340 30254 3352
rect 30653 3349 30665 3352
rect 30699 3349 30711 3383
rect 30653 3343 30711 3349
rect 1104 3290 34316 3312
rect 1104 3238 6517 3290
rect 6569 3238 6581 3290
rect 6633 3238 6645 3290
rect 6697 3238 6709 3290
rect 6761 3238 17588 3290
rect 17640 3238 17652 3290
rect 17704 3238 17716 3290
rect 17768 3238 17780 3290
rect 17832 3238 28658 3290
rect 28710 3238 28722 3290
rect 28774 3238 28786 3290
rect 28838 3238 28850 3290
rect 28902 3238 34316 3290
rect 1104 3216 34316 3238
rect 17402 3136 17408 3188
rect 17460 3176 17466 3188
rect 17497 3179 17555 3185
rect 17497 3176 17509 3179
rect 17460 3148 17509 3176
rect 17460 3136 17466 3148
rect 17497 3145 17509 3148
rect 17543 3145 17555 3179
rect 19150 3176 19156 3188
rect 17497 3139 17555 3145
rect 18064 3148 19156 3176
rect 18064 3108 18092 3148
rect 19150 3136 19156 3148
rect 19208 3176 19214 3188
rect 20533 3179 20591 3185
rect 20533 3176 20545 3179
rect 19208 3148 20545 3176
rect 19208 3136 19214 3148
rect 20533 3145 20545 3148
rect 20579 3145 20591 3179
rect 20533 3139 20591 3145
rect 26510 3136 26516 3188
rect 26568 3176 26574 3188
rect 30193 3179 30251 3185
rect 26568 3148 29776 3176
rect 26568 3136 26574 3148
rect 17420 3080 18092 3108
rect 17420 3049 17448 3080
rect 17405 3043 17463 3049
rect 17405 3009 17417 3043
rect 17451 3009 17463 3043
rect 17586 3040 17592 3052
rect 17547 3012 17592 3040
rect 17405 3003 17463 3009
rect 17586 3000 17592 3012
rect 17644 3000 17650 3052
rect 28460 3049 28488 3148
rect 29748 3108 29776 3148
rect 30193 3145 30205 3179
rect 30239 3176 30251 3179
rect 30282 3176 30288 3188
rect 30239 3148 30288 3176
rect 30239 3145 30251 3148
rect 30193 3139 30251 3145
rect 30282 3136 30288 3148
rect 30340 3136 30346 3188
rect 30745 3179 30803 3185
rect 30745 3145 30757 3179
rect 30791 3176 30803 3179
rect 31202 3176 31208 3188
rect 30791 3148 31208 3176
rect 30791 3145 30803 3148
rect 30745 3139 30803 3145
rect 31202 3136 31208 3148
rect 31260 3136 31266 3188
rect 31570 3108 31576 3120
rect 29748 3080 31576 3108
rect 31570 3068 31576 3080
rect 31628 3068 31634 3120
rect 20717 3043 20775 3049
rect 20717 3009 20729 3043
rect 20763 3040 20775 3043
rect 21269 3043 21327 3049
rect 21269 3040 21281 3043
rect 20763 3012 21281 3040
rect 20763 3009 20775 3012
rect 20717 3003 20775 3009
rect 21269 3009 21281 3012
rect 21315 3009 21327 3043
rect 21269 3003 21327 3009
rect 28445 3043 28503 3049
rect 28445 3009 28457 3043
rect 28491 3009 28503 3043
rect 28445 3003 28503 3009
rect 28721 3043 28779 3049
rect 28721 3009 28733 3043
rect 28767 3040 28779 3043
rect 29086 3040 29092 3052
rect 28767 3012 29092 3040
rect 28767 3009 28779 3012
rect 28721 3003 28779 3009
rect 29086 3000 29092 3012
rect 29144 3000 29150 3052
rect 17218 2932 17224 2984
rect 17276 2972 17282 2984
rect 18322 2981 18328 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 17276 2944 17325 2972
rect 17276 2932 17282 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 18049 2975 18107 2981
rect 18049 2941 18061 2975
rect 18095 2941 18107 2975
rect 18316 2972 18328 2981
rect 18283 2944 18328 2972
rect 18049 2935 18107 2941
rect 18316 2935 18328 2944
rect 17126 2864 17132 2916
rect 17184 2904 17190 2916
rect 18064 2904 18092 2935
rect 18322 2932 18328 2935
rect 18380 2932 18386 2984
rect 20438 2972 20444 2984
rect 20399 2944 20444 2972
rect 20438 2932 20444 2944
rect 20496 2932 20502 2984
rect 21177 2975 21235 2981
rect 21177 2941 21189 2975
rect 21223 2941 21235 2975
rect 21177 2935 21235 2941
rect 21361 2975 21419 2981
rect 21361 2941 21373 2975
rect 21407 2972 21419 2975
rect 21910 2972 21916 2984
rect 21407 2944 21916 2972
rect 21407 2941 21419 2944
rect 21361 2935 21419 2941
rect 17184 2876 19840 2904
rect 17184 2864 17190 2876
rect 19426 2836 19432 2848
rect 19387 2808 19432 2836
rect 19426 2796 19432 2808
rect 19484 2796 19490 2848
rect 19812 2836 19840 2876
rect 19886 2864 19892 2916
rect 19944 2904 19950 2916
rect 21192 2904 21220 2935
rect 21910 2932 21916 2944
rect 21968 2932 21974 2984
rect 30650 2972 30656 2984
rect 30611 2944 30656 2972
rect 30650 2932 30656 2944
rect 30708 2932 30714 2984
rect 32858 2904 32864 2916
rect 19944 2876 21220 2904
rect 29946 2890 32864 2904
rect 29932 2876 32864 2890
rect 19944 2864 19950 2876
rect 20530 2836 20536 2848
rect 19812 2808 20536 2836
rect 20530 2796 20536 2808
rect 20588 2796 20594 2848
rect 20714 2836 20720 2848
rect 20675 2808 20720 2836
rect 20714 2796 20720 2808
rect 20772 2796 20778 2848
rect 27522 2796 27528 2848
rect 27580 2836 27586 2848
rect 29932 2836 29960 2876
rect 32858 2864 32864 2876
rect 32916 2864 32922 2916
rect 27580 2808 29960 2836
rect 27580 2796 27586 2808
rect 1104 2746 34316 2768
rect 1104 2694 12052 2746
rect 12104 2694 12116 2746
rect 12168 2694 12180 2746
rect 12232 2694 12244 2746
rect 12296 2694 23123 2746
rect 23175 2694 23187 2746
rect 23239 2694 23251 2746
rect 23303 2694 23315 2746
rect 23367 2694 34316 2746
rect 1104 2672 34316 2694
rect 5718 2632 5724 2644
rect 5679 2604 5724 2632
rect 5718 2592 5724 2604
rect 5776 2592 5782 2644
rect 6886 2604 11468 2632
rect 1949 2567 2007 2573
rect 1949 2533 1961 2567
rect 1995 2564 2007 2567
rect 6886 2564 6914 2604
rect 11238 2564 11244 2576
rect 1995 2536 6914 2564
rect 11199 2536 11244 2564
rect 1995 2533 2007 2536
rect 1949 2527 2007 2533
rect 11238 2524 11244 2536
rect 11296 2524 11302 2576
rect 11440 2564 11468 2604
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 13817 2635 13875 2641
rect 13817 2632 13829 2635
rect 12492 2604 13829 2632
rect 12492 2592 12498 2604
rect 13817 2601 13829 2604
rect 13863 2601 13875 2635
rect 13817 2595 13875 2601
rect 17586 2592 17592 2644
rect 17644 2632 17650 2644
rect 17681 2635 17739 2641
rect 17681 2632 17693 2635
rect 17644 2604 17693 2632
rect 17644 2592 17650 2604
rect 17681 2601 17693 2604
rect 17727 2601 17739 2635
rect 18414 2632 18420 2644
rect 18375 2604 18420 2632
rect 17681 2595 17739 2601
rect 18414 2592 18420 2604
rect 18472 2592 18478 2644
rect 21910 2632 21916 2644
rect 21871 2604 21916 2632
rect 21910 2592 21916 2604
rect 21968 2632 21974 2644
rect 21968 2604 23152 2632
rect 21968 2592 21974 2604
rect 16022 2564 16028 2576
rect 11440 2536 16028 2564
rect 16022 2524 16028 2536
rect 16080 2524 16086 2576
rect 16482 2564 16488 2576
rect 16443 2536 16488 2564
rect 16482 2524 16488 2536
rect 16540 2524 16546 2576
rect 19153 2567 19211 2573
rect 19153 2533 19165 2567
rect 19199 2564 19211 2567
rect 19426 2564 19432 2576
rect 19199 2536 19432 2564
rect 19199 2533 19211 2536
rect 19153 2527 19211 2533
rect 2774 2456 2780 2508
rect 2832 2496 2838 2508
rect 2869 2499 2927 2505
rect 2869 2496 2881 2499
rect 2832 2468 2881 2496
rect 2832 2456 2838 2468
rect 2869 2465 2881 2468
rect 2915 2465 2927 2499
rect 5534 2496 5540 2508
rect 5495 2468 5540 2496
rect 2869 2459 2927 2465
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 8481 2499 8539 2505
rect 8481 2465 8493 2499
rect 8527 2465 8539 2499
rect 8481 2459 8539 2465
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 8496 2428 8524 2459
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 14001 2499 14059 2505
rect 14001 2496 14013 2499
rect 13872 2468 14013 2496
rect 13872 2456 13878 2468
rect 14001 2465 14013 2468
rect 14047 2465 14059 2499
rect 17589 2499 17647 2505
rect 17589 2496 17601 2499
rect 14001 2459 14059 2465
rect 16546 2468 17601 2496
rect 16114 2428 16120 2440
rect 3099 2400 6914 2428
rect 8496 2400 16120 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 474 2320 480 2372
rect 532 2360 538 2372
rect 1765 2363 1823 2369
rect 1765 2360 1777 2363
rect 532 2332 1777 2360
rect 532 2320 538 2332
rect 1765 2329 1777 2332
rect 1811 2329 1823 2363
rect 1765 2323 1823 2329
rect 6886 2292 6914 2400
rect 16114 2388 16120 2400
rect 16172 2428 16178 2440
rect 16546 2428 16574 2468
rect 17589 2465 17601 2468
rect 17635 2465 17647 2499
rect 17589 2459 17647 2465
rect 17773 2499 17831 2505
rect 17773 2465 17785 2499
rect 17819 2496 17831 2499
rect 18417 2499 18475 2505
rect 18417 2496 18429 2499
rect 17819 2468 18429 2496
rect 17819 2465 17831 2468
rect 17773 2459 17831 2465
rect 18417 2465 18429 2468
rect 18463 2465 18475 2499
rect 18417 2459 18475 2465
rect 18601 2499 18659 2505
rect 18601 2465 18613 2499
rect 18647 2496 18659 2499
rect 19168 2496 19196 2527
rect 19426 2524 19432 2536
rect 19484 2524 19490 2576
rect 20714 2524 20720 2576
rect 20772 2573 20778 2576
rect 23124 2573 23152 2604
rect 20772 2567 20836 2573
rect 20772 2533 20790 2567
rect 20824 2533 20836 2567
rect 20772 2527 20836 2533
rect 23109 2567 23167 2573
rect 23109 2533 23121 2567
rect 23155 2533 23167 2567
rect 25774 2564 25780 2576
rect 25735 2536 25780 2564
rect 23109 2527 23167 2533
rect 20772 2524 20778 2527
rect 25774 2524 25780 2536
rect 25832 2524 25838 2576
rect 28442 2564 28448 2576
rect 28403 2536 28448 2564
rect 28442 2524 28448 2536
rect 28500 2524 28506 2576
rect 30374 2524 30380 2576
rect 30432 2564 30438 2576
rect 31113 2567 31171 2573
rect 31113 2564 31125 2567
rect 30432 2536 31125 2564
rect 30432 2524 30438 2536
rect 31113 2533 31125 2536
rect 31159 2533 31171 2567
rect 31754 2564 31760 2576
rect 31715 2536 31760 2564
rect 31113 2527 31171 2533
rect 31754 2524 31760 2536
rect 31812 2524 31818 2576
rect 32490 2564 32496 2576
rect 32451 2536 32496 2564
rect 32490 2524 32496 2536
rect 32548 2524 32554 2576
rect 20530 2496 20536 2508
rect 18647 2468 19196 2496
rect 20491 2468 20536 2496
rect 18647 2465 18659 2468
rect 18601 2459 18659 2465
rect 16172 2400 16574 2428
rect 18432 2428 18460 2459
rect 20530 2456 20536 2468
rect 20588 2456 20594 2508
rect 19978 2428 19984 2440
rect 18432 2400 19984 2428
rect 16172 2388 16178 2400
rect 19978 2388 19984 2400
rect 20036 2388 20042 2440
rect 8294 2360 8300 2372
rect 8255 2332 8300 2360
rect 8294 2320 8300 2332
rect 8352 2320 8358 2372
rect 11054 2360 11060 2372
rect 11015 2332 11060 2360
rect 11054 2320 11060 2332
rect 11112 2320 11118 2372
rect 19334 2360 19340 2372
rect 19295 2332 19340 2360
rect 19334 2320 19340 2332
rect 19392 2320 19398 2372
rect 22094 2320 22100 2372
rect 22152 2360 22158 2372
rect 22925 2363 22983 2369
rect 22925 2360 22937 2363
rect 22152 2332 22937 2360
rect 22152 2320 22158 2332
rect 22925 2329 22937 2332
rect 22971 2329 22983 2363
rect 22925 2323 22983 2329
rect 24854 2320 24860 2372
rect 24912 2360 24918 2372
rect 25593 2363 25651 2369
rect 25593 2360 25605 2363
rect 24912 2332 25605 2360
rect 24912 2320 24918 2332
rect 25593 2329 25605 2332
rect 25639 2329 25651 2363
rect 25593 2323 25651 2329
rect 27614 2320 27620 2372
rect 27672 2360 27678 2372
rect 28261 2363 28319 2369
rect 28261 2360 28273 2363
rect 27672 2332 28273 2360
rect 27672 2320 27678 2332
rect 28261 2329 28273 2332
rect 28307 2329 28319 2363
rect 28261 2323 28319 2329
rect 30374 2320 30380 2372
rect 30432 2360 30438 2372
rect 30929 2363 30987 2369
rect 30929 2360 30941 2363
rect 30432 2332 30941 2360
rect 30432 2320 30438 2332
rect 30929 2329 30941 2332
rect 30975 2329 30987 2363
rect 31938 2360 31944 2372
rect 31899 2332 31944 2360
rect 30929 2323 30987 2329
rect 31938 2320 31944 2332
rect 31996 2320 32002 2372
rect 32674 2360 32680 2372
rect 32635 2332 32680 2360
rect 32674 2320 32680 2332
rect 32732 2320 32738 2372
rect 16298 2292 16304 2304
rect 6886 2264 16304 2292
rect 16298 2252 16304 2264
rect 16356 2252 16362 2304
rect 16574 2252 16580 2304
rect 16632 2292 16638 2304
rect 16632 2264 16677 2292
rect 16632 2252 16638 2264
rect 1104 2202 34316 2224
rect 1104 2150 6517 2202
rect 6569 2150 6581 2202
rect 6633 2150 6645 2202
rect 6697 2150 6709 2202
rect 6761 2150 17588 2202
rect 17640 2150 17652 2202
rect 17704 2150 17716 2202
rect 17768 2150 17780 2202
rect 17832 2150 28658 2202
rect 28710 2150 28722 2202
rect 28774 2150 28786 2202
rect 28838 2150 28850 2202
rect 28902 2150 34316 2202
rect 1104 2128 34316 2150
<< via1 >>
rect 7104 35436 7156 35488
rect 15844 35436 15896 35488
rect 12052 35334 12104 35386
rect 12116 35334 12168 35386
rect 12180 35334 12232 35386
rect 12244 35334 12296 35386
rect 23123 35334 23175 35386
rect 23187 35334 23239 35386
rect 23251 35334 23303 35386
rect 23315 35334 23367 35386
rect 7104 35232 7156 35284
rect 12624 35232 12676 35284
rect 21640 35232 21692 35284
rect 24400 35232 24452 35284
rect 10600 35207 10652 35216
rect 1400 35139 1452 35148
rect 1400 35105 1409 35139
rect 1409 35105 1443 35139
rect 1443 35105 1452 35139
rect 1400 35096 1452 35105
rect 2780 35139 2832 35148
rect 2780 35105 2789 35139
rect 2789 35105 2823 35139
rect 2823 35105 2832 35139
rect 2780 35096 2832 35105
rect 5080 35139 5132 35148
rect 5080 35105 5089 35139
rect 5089 35105 5123 35139
rect 5123 35105 5132 35139
rect 5080 35096 5132 35105
rect 7840 35096 7892 35148
rect 8392 35096 8444 35148
rect 2964 34935 3016 34944
rect 2964 34901 2973 34935
rect 2973 34901 3007 34935
rect 3007 34901 3016 34935
rect 2964 34892 3016 34901
rect 8208 34960 8260 35012
rect 10600 35173 10609 35207
rect 10609 35173 10643 35207
rect 10643 35173 10652 35207
rect 10600 35164 10652 35173
rect 13360 35207 13412 35216
rect 13360 35173 13369 35207
rect 13369 35173 13403 35207
rect 13403 35173 13412 35207
rect 13360 35164 13412 35173
rect 13452 35164 13504 35216
rect 27068 35164 27120 35216
rect 27160 35164 27212 35216
rect 32680 35164 32732 35216
rect 14464 35096 14516 35148
rect 16120 35096 16172 35148
rect 18880 35139 18932 35148
rect 18880 35105 18889 35139
rect 18889 35105 18923 35139
rect 18923 35105 18932 35139
rect 18880 35096 18932 35105
rect 21824 35139 21876 35148
rect 21824 35105 21833 35139
rect 21833 35105 21867 35139
rect 21867 35105 21876 35139
rect 21824 35096 21876 35105
rect 14280 35028 14332 35080
rect 20076 35028 20128 35080
rect 29920 35096 29972 35148
rect 34980 35096 35032 35148
rect 29276 35028 29328 35080
rect 12532 34960 12584 35012
rect 8484 34892 8536 34944
rect 8668 34892 8720 34944
rect 15292 34892 15344 34944
rect 18880 34892 18932 34944
rect 29460 34892 29512 34944
rect 32312 34892 32364 34944
rect 32496 34935 32548 34944
rect 32496 34901 32505 34935
rect 32505 34901 32539 34935
rect 32539 34901 32548 34935
rect 32496 34892 32548 34901
rect 6517 34790 6569 34842
rect 6581 34790 6633 34842
rect 6645 34790 6697 34842
rect 6709 34790 6761 34842
rect 17588 34790 17640 34842
rect 17652 34790 17704 34842
rect 17716 34790 17768 34842
rect 17780 34790 17832 34842
rect 28658 34790 28710 34842
rect 28722 34790 28774 34842
rect 28786 34790 28838 34842
rect 28850 34790 28902 34842
rect 8392 34731 8444 34740
rect 8392 34697 8401 34731
rect 8401 34697 8435 34731
rect 8435 34697 8444 34731
rect 8392 34688 8444 34697
rect 8484 34688 8536 34740
rect 2964 34620 3016 34672
rect 7196 34552 7248 34604
rect 9680 34620 9732 34672
rect 12532 34552 12584 34604
rect 27068 34688 27120 34740
rect 16396 34620 16448 34672
rect 9956 34527 10008 34536
rect 9956 34493 9965 34527
rect 9965 34493 9999 34527
rect 9999 34493 10008 34527
rect 9956 34484 10008 34493
rect 10508 34484 10560 34536
rect 12992 34484 13044 34536
rect 13820 34527 13872 34536
rect 13820 34493 13829 34527
rect 13829 34493 13863 34527
rect 13863 34493 13872 34527
rect 13820 34484 13872 34493
rect 19892 34552 19944 34604
rect 17132 34484 17184 34536
rect 19432 34527 19484 34536
rect 19432 34493 19441 34527
rect 19441 34493 19475 34527
rect 19475 34493 19484 34527
rect 19432 34484 19484 34493
rect 23020 34527 23072 34536
rect 8208 34348 8260 34400
rect 10140 34391 10192 34400
rect 10140 34357 10149 34391
rect 10149 34357 10183 34391
rect 10183 34357 10192 34391
rect 10140 34348 10192 34357
rect 12440 34391 12492 34400
rect 12440 34357 12449 34391
rect 12449 34357 12483 34391
rect 12483 34357 12492 34391
rect 12440 34348 12492 34357
rect 12532 34391 12584 34400
rect 12532 34357 12541 34391
rect 12541 34357 12575 34391
rect 12575 34357 12584 34391
rect 20996 34416 21048 34468
rect 23020 34493 23029 34527
rect 23029 34493 23063 34527
rect 23063 34493 23072 34527
rect 23020 34484 23072 34493
rect 29460 34527 29512 34536
rect 29460 34493 29469 34527
rect 29469 34493 29503 34527
rect 29503 34493 29512 34527
rect 29460 34484 29512 34493
rect 12532 34348 12584 34357
rect 20720 34348 20772 34400
rect 21916 34348 21968 34400
rect 23756 34348 23808 34400
rect 12052 34246 12104 34298
rect 12116 34246 12168 34298
rect 12180 34246 12232 34298
rect 12244 34246 12296 34298
rect 23123 34246 23175 34298
rect 23187 34246 23239 34298
rect 23251 34246 23303 34298
rect 23315 34246 23367 34298
rect 12440 34144 12492 34196
rect 12532 34144 12584 34196
rect 13452 34144 13504 34196
rect 23020 34144 23072 34196
rect 23756 34187 23808 34196
rect 23756 34153 23765 34187
rect 23765 34153 23799 34187
rect 23799 34153 23808 34187
rect 23756 34144 23808 34153
rect 10140 34119 10192 34128
rect 10140 34085 10174 34119
rect 10174 34085 10192 34119
rect 10140 34076 10192 34085
rect 13452 34051 13504 34060
rect 13452 34017 13461 34051
rect 13461 34017 13495 34051
rect 13495 34017 13504 34051
rect 13452 34008 13504 34017
rect 13820 34008 13872 34060
rect 16304 34008 16356 34060
rect 17132 34051 17184 34060
rect 17132 34017 17141 34051
rect 17141 34017 17175 34051
rect 17175 34017 17184 34051
rect 17132 34008 17184 34017
rect 9680 33940 9732 33992
rect 12808 33983 12860 33992
rect 12808 33949 12817 33983
rect 12817 33949 12851 33983
rect 12851 33949 12860 33983
rect 12808 33940 12860 33949
rect 18052 33940 18104 33992
rect 11244 33847 11296 33856
rect 11244 33813 11253 33847
rect 11253 33813 11287 33847
rect 11287 33813 11296 33847
rect 11244 33804 11296 33813
rect 13544 33847 13596 33856
rect 13544 33813 13553 33847
rect 13553 33813 13587 33847
rect 13587 33813 13596 33847
rect 13544 33804 13596 33813
rect 17960 33804 18012 33856
rect 20720 34076 20772 34128
rect 21916 34076 21968 34128
rect 23572 34008 23624 34060
rect 20996 33983 21048 33992
rect 20996 33949 21005 33983
rect 21005 33949 21039 33983
rect 21039 33949 21048 33983
rect 20996 33940 21048 33949
rect 21640 33940 21692 33992
rect 23940 33983 23992 33992
rect 23940 33949 23949 33983
rect 23949 33949 23983 33983
rect 23983 33949 23992 33983
rect 23940 33940 23992 33949
rect 19340 33804 19392 33856
rect 21180 33804 21232 33856
rect 23572 33804 23624 33856
rect 6517 33702 6569 33754
rect 6581 33702 6633 33754
rect 6645 33702 6697 33754
rect 6709 33702 6761 33754
rect 17588 33702 17640 33754
rect 17652 33702 17704 33754
rect 17716 33702 17768 33754
rect 17780 33702 17832 33754
rect 28658 33702 28710 33754
rect 28722 33702 28774 33754
rect 28786 33702 28838 33754
rect 28850 33702 28902 33754
rect 8208 33643 8260 33652
rect 8208 33609 8217 33643
rect 8217 33609 8251 33643
rect 8251 33609 8260 33643
rect 8208 33600 8260 33609
rect 12532 33600 12584 33652
rect 18052 33600 18104 33652
rect 19432 33643 19484 33652
rect 19432 33609 19441 33643
rect 19441 33609 19475 33643
rect 19475 33609 19484 33643
rect 19432 33600 19484 33609
rect 21640 33643 21692 33652
rect 21640 33609 21649 33643
rect 21649 33609 21683 33643
rect 21683 33609 21692 33643
rect 21640 33600 21692 33609
rect 21824 33532 21876 33584
rect 5080 33464 5132 33516
rect 2964 33396 3016 33448
rect 3976 33439 4028 33448
rect 3056 33328 3108 33380
rect 3976 33405 3985 33439
rect 3985 33405 4019 33439
rect 4019 33405 4028 33439
rect 3976 33396 4028 33405
rect 8668 33439 8720 33448
rect 8668 33405 8677 33439
rect 8677 33405 8711 33439
rect 8711 33405 8720 33439
rect 8668 33396 8720 33405
rect 8944 33439 8996 33448
rect 8944 33405 8953 33439
rect 8953 33405 8987 33439
rect 8987 33405 8996 33439
rect 8944 33396 8996 33405
rect 9496 33439 9548 33448
rect 9496 33405 9505 33439
rect 9505 33405 9539 33439
rect 9539 33405 9548 33439
rect 9496 33396 9548 33405
rect 10416 33396 10468 33448
rect 13544 33464 13596 33516
rect 13820 33464 13872 33516
rect 19892 33507 19944 33516
rect 12532 33396 12584 33448
rect 13268 33439 13320 33448
rect 13268 33405 13277 33439
rect 13277 33405 13311 33439
rect 13311 33405 13320 33439
rect 13268 33396 13320 33405
rect 13452 33439 13504 33448
rect 13452 33405 13461 33439
rect 13461 33405 13495 33439
rect 13495 33405 13504 33439
rect 13452 33396 13504 33405
rect 18604 33396 18656 33448
rect 19892 33473 19901 33507
rect 19901 33473 19935 33507
rect 19935 33473 19944 33507
rect 19892 33464 19944 33473
rect 20720 33464 20772 33516
rect 21180 33507 21232 33516
rect 21180 33473 21189 33507
rect 21189 33473 21223 33507
rect 21223 33473 21232 33507
rect 21180 33464 21232 33473
rect 25320 33439 25372 33448
rect 25320 33405 25329 33439
rect 25329 33405 25363 33439
rect 25363 33405 25372 33439
rect 25320 33396 25372 33405
rect 27804 33396 27856 33448
rect 29276 33396 29328 33448
rect 33600 33439 33652 33448
rect 33600 33405 33609 33439
rect 33609 33405 33643 33439
rect 33643 33405 33652 33439
rect 33600 33396 33652 33405
rect 5448 33328 5500 33380
rect 9956 33328 10008 33380
rect 3608 33260 3660 33312
rect 6920 33260 6972 33312
rect 7748 33303 7800 33312
rect 7748 33269 7757 33303
rect 7757 33269 7791 33303
rect 7791 33269 7800 33303
rect 7748 33260 7800 33269
rect 8576 33260 8628 33312
rect 8760 33303 8812 33312
rect 8760 33269 8769 33303
rect 8769 33269 8803 33303
rect 8803 33269 8812 33303
rect 8760 33260 8812 33269
rect 11244 33260 11296 33312
rect 14740 33328 14792 33380
rect 21916 33328 21968 33380
rect 24308 33328 24360 33380
rect 28172 33371 28224 33380
rect 28172 33337 28181 33371
rect 28181 33337 28215 33371
rect 28215 33337 28224 33371
rect 28172 33328 28224 33337
rect 30012 33328 30064 33380
rect 15476 33260 15528 33312
rect 18512 33303 18564 33312
rect 18512 33269 18521 33303
rect 18521 33269 18555 33303
rect 18555 33269 18564 33303
rect 18512 33260 18564 33269
rect 19340 33260 19392 33312
rect 19800 33303 19852 33312
rect 19800 33269 19809 33303
rect 19809 33269 19843 33303
rect 19843 33269 19852 33303
rect 19800 33260 19852 33269
rect 21272 33303 21324 33312
rect 21272 33269 21281 33303
rect 21281 33269 21315 33303
rect 21315 33269 21324 33303
rect 21272 33260 21324 33269
rect 23664 33260 23716 33312
rect 33416 33303 33468 33312
rect 33416 33269 33425 33303
rect 33425 33269 33459 33303
rect 33459 33269 33468 33303
rect 33416 33260 33468 33269
rect 12052 33158 12104 33210
rect 12116 33158 12168 33210
rect 12180 33158 12232 33210
rect 12244 33158 12296 33210
rect 23123 33158 23175 33210
rect 23187 33158 23239 33210
rect 23251 33158 23303 33210
rect 23315 33158 23367 33210
rect 7656 33056 7708 33108
rect 7748 33056 7800 33108
rect 10508 33099 10560 33108
rect 10508 33065 10517 33099
rect 10517 33065 10551 33099
rect 10551 33065 10560 33099
rect 10508 33056 10560 33065
rect 3884 32988 3936 33040
rect 17408 33056 17460 33108
rect 1400 32963 1452 32972
rect 1400 32929 1409 32963
rect 1409 32929 1443 32963
rect 1443 32929 1452 32963
rect 1400 32920 1452 32929
rect 5632 32963 5684 32972
rect 5632 32929 5650 32963
rect 5650 32929 5684 32963
rect 5632 32920 5684 32929
rect 8300 32920 8352 32972
rect 17776 32988 17828 33040
rect 18512 32988 18564 33040
rect 23572 33031 23624 33040
rect 23572 32997 23581 33031
rect 23581 32997 23615 33031
rect 23615 32997 23624 33031
rect 23572 32988 23624 32997
rect 10232 32920 10284 32972
rect 10416 32920 10468 32972
rect 4528 32759 4580 32768
rect 4528 32725 4537 32759
rect 4537 32725 4571 32759
rect 4571 32725 4580 32759
rect 4528 32716 4580 32725
rect 6920 32716 6972 32768
rect 9680 32852 9732 32904
rect 9956 32852 10008 32904
rect 10324 32852 10376 32904
rect 11244 32920 11296 32972
rect 13544 32920 13596 32972
rect 14832 32920 14884 32972
rect 16304 32920 16356 32972
rect 23756 32920 23808 32972
rect 33416 32963 33468 32972
rect 33416 32929 33425 32963
rect 33425 32929 33459 32963
rect 33459 32929 33468 32963
rect 33416 32920 33468 32929
rect 12900 32895 12952 32904
rect 12900 32861 12909 32895
rect 12909 32861 12943 32895
rect 12943 32861 12952 32895
rect 12900 32852 12952 32861
rect 12992 32895 13044 32904
rect 12992 32861 13001 32895
rect 13001 32861 13035 32895
rect 13035 32861 13044 32895
rect 15200 32895 15252 32904
rect 12992 32852 13044 32861
rect 15200 32861 15209 32895
rect 15209 32861 15243 32895
rect 15243 32861 15252 32895
rect 15200 32852 15252 32861
rect 17960 32852 18012 32904
rect 19800 32852 19852 32904
rect 21272 32852 21324 32904
rect 22836 32852 22888 32904
rect 19156 32784 19208 32836
rect 23664 32784 23716 32836
rect 8484 32759 8536 32768
rect 8484 32725 8493 32759
rect 8493 32725 8527 32759
rect 8527 32725 8536 32759
rect 8484 32716 8536 32725
rect 8944 32716 8996 32768
rect 9588 32716 9640 32768
rect 10048 32716 10100 32768
rect 14188 32716 14240 32768
rect 19892 32716 19944 32768
rect 20260 32759 20312 32768
rect 20260 32725 20269 32759
rect 20269 32725 20303 32759
rect 20303 32725 20312 32759
rect 20260 32716 20312 32725
rect 20444 32759 20496 32768
rect 20444 32725 20453 32759
rect 20453 32725 20487 32759
rect 20487 32725 20496 32759
rect 20444 32716 20496 32725
rect 33508 32759 33560 32768
rect 33508 32725 33517 32759
rect 33517 32725 33551 32759
rect 33551 32725 33560 32759
rect 33508 32716 33560 32725
rect 6517 32614 6569 32666
rect 6581 32614 6633 32666
rect 6645 32614 6697 32666
rect 6709 32614 6761 32666
rect 17588 32614 17640 32666
rect 17652 32614 17704 32666
rect 17716 32614 17768 32666
rect 17780 32614 17832 32666
rect 28658 32614 28710 32666
rect 28722 32614 28774 32666
rect 28786 32614 28838 32666
rect 28850 32614 28902 32666
rect 5080 32555 5132 32564
rect 5080 32521 5089 32555
rect 5089 32521 5123 32555
rect 5123 32521 5132 32555
rect 5080 32512 5132 32521
rect 8300 32555 8352 32564
rect 8300 32521 8309 32555
rect 8309 32521 8343 32555
rect 8343 32521 8352 32555
rect 8300 32512 8352 32521
rect 8576 32512 8628 32564
rect 12900 32512 12952 32564
rect 13544 32555 13596 32564
rect 5356 32376 5408 32428
rect 7472 32419 7524 32428
rect 7472 32385 7481 32419
rect 7481 32385 7515 32419
rect 7515 32385 7524 32419
rect 7472 32376 7524 32385
rect 12532 32419 12584 32428
rect 3608 32351 3660 32360
rect 3608 32317 3626 32351
rect 3626 32317 3660 32351
rect 3884 32351 3936 32360
rect 3608 32308 3660 32317
rect 3884 32317 3893 32351
rect 3893 32317 3927 32351
rect 3927 32317 3936 32351
rect 3884 32308 3936 32317
rect 6920 32308 6972 32360
rect 8484 32351 8536 32360
rect 8484 32317 8493 32351
rect 8493 32317 8527 32351
rect 8527 32317 8536 32351
rect 8484 32308 8536 32317
rect 12532 32385 12541 32419
rect 12541 32385 12575 32419
rect 12575 32385 12584 32419
rect 12532 32376 12584 32385
rect 8760 32240 8812 32292
rect 9588 32308 9640 32360
rect 9680 32308 9732 32360
rect 10048 32351 10100 32360
rect 10048 32317 10082 32351
rect 10082 32317 10100 32351
rect 10048 32308 10100 32317
rect 13544 32521 13553 32555
rect 13553 32521 13587 32555
rect 13587 32521 13596 32555
rect 13544 32512 13596 32521
rect 14832 32555 14884 32564
rect 14832 32521 14841 32555
rect 14841 32521 14875 32555
rect 14875 32521 14884 32555
rect 14832 32512 14884 32521
rect 33508 32512 33560 32564
rect 17960 32487 18012 32496
rect 17960 32453 17969 32487
rect 17969 32453 18003 32487
rect 18003 32453 18012 32487
rect 17960 32444 18012 32453
rect 19340 32487 19392 32496
rect 19340 32453 19349 32487
rect 19349 32453 19383 32487
rect 19383 32453 19392 32487
rect 19340 32444 19392 32453
rect 21272 32444 21324 32496
rect 25320 32444 25372 32496
rect 28172 32444 28224 32496
rect 15292 32419 15344 32428
rect 15292 32385 15301 32419
rect 15301 32385 15335 32419
rect 15335 32385 15344 32419
rect 15292 32376 15344 32385
rect 15200 32351 15252 32360
rect 9956 32240 10008 32292
rect 3148 32172 3200 32224
rect 4528 32172 4580 32224
rect 5540 32215 5592 32224
rect 5540 32181 5549 32215
rect 5549 32181 5583 32215
rect 5583 32181 5592 32215
rect 5540 32172 5592 32181
rect 5724 32172 5776 32224
rect 7288 32215 7340 32224
rect 7288 32181 7297 32215
rect 7297 32181 7331 32215
rect 7331 32181 7340 32215
rect 7288 32172 7340 32181
rect 7380 32215 7432 32224
rect 7380 32181 7389 32215
rect 7389 32181 7423 32215
rect 7423 32181 7432 32215
rect 7380 32172 7432 32181
rect 9588 32172 9640 32224
rect 13268 32240 13320 32292
rect 15200 32317 15209 32351
rect 15209 32317 15243 32351
rect 15243 32317 15252 32351
rect 15200 32308 15252 32317
rect 18144 32376 18196 32428
rect 18604 32419 18656 32428
rect 18604 32385 18613 32419
rect 18613 32385 18647 32419
rect 18647 32385 18656 32419
rect 18604 32376 18656 32385
rect 19156 32351 19208 32360
rect 19156 32317 19165 32351
rect 19165 32317 19199 32351
rect 19199 32317 19208 32351
rect 19156 32308 19208 32317
rect 20444 32376 20496 32428
rect 23480 32376 23532 32428
rect 23940 32376 23992 32428
rect 26608 32376 26660 32428
rect 29460 32419 29512 32428
rect 29460 32385 29469 32419
rect 29469 32385 29503 32419
rect 29503 32385 29512 32419
rect 29460 32376 29512 32385
rect 20168 32351 20220 32360
rect 11152 32215 11204 32224
rect 11152 32181 11161 32215
rect 11161 32181 11195 32215
rect 11195 32181 11204 32215
rect 11152 32172 11204 32181
rect 12440 32172 12492 32224
rect 12992 32172 13044 32224
rect 13176 32172 13228 32224
rect 18512 32240 18564 32292
rect 17960 32172 18012 32224
rect 20168 32317 20177 32351
rect 20177 32317 20211 32351
rect 20211 32317 20220 32351
rect 20168 32308 20220 32317
rect 23664 32308 23716 32360
rect 27804 32308 27856 32360
rect 21180 32240 21232 32292
rect 21916 32240 21968 32292
rect 23756 32240 23808 32292
rect 26700 32240 26752 32292
rect 30472 32240 30524 32292
rect 30656 32240 30708 32292
rect 20996 32172 21048 32224
rect 21364 32172 21416 32224
rect 22100 32172 22152 32224
rect 22836 32215 22888 32224
rect 22836 32181 22845 32215
rect 22845 32181 22879 32215
rect 22879 32181 22888 32215
rect 22836 32172 22888 32181
rect 23020 32172 23072 32224
rect 25872 32215 25924 32224
rect 25872 32181 25881 32215
rect 25881 32181 25915 32215
rect 25915 32181 25924 32215
rect 25872 32172 25924 32181
rect 26240 32215 26292 32224
rect 26240 32181 26249 32215
rect 26249 32181 26283 32215
rect 26283 32181 26292 32215
rect 29276 32215 29328 32224
rect 26240 32172 26292 32181
rect 29276 32181 29285 32215
rect 29285 32181 29319 32215
rect 29319 32181 29328 32215
rect 29276 32172 29328 32181
rect 30748 32172 30800 32224
rect 12052 32070 12104 32122
rect 12116 32070 12168 32122
rect 12180 32070 12232 32122
rect 12244 32070 12296 32122
rect 23123 32070 23175 32122
rect 23187 32070 23239 32122
rect 23251 32070 23303 32122
rect 23315 32070 23367 32122
rect 3976 31968 4028 32020
rect 5632 31968 5684 32020
rect 7380 31968 7432 32020
rect 9588 32011 9640 32020
rect 9588 31977 9597 32011
rect 9597 31977 9631 32011
rect 9631 31977 9640 32011
rect 9588 31968 9640 31977
rect 10232 32011 10284 32020
rect 10232 31977 10241 32011
rect 10241 31977 10275 32011
rect 10275 31977 10284 32011
rect 10232 31968 10284 31977
rect 12440 32011 12492 32020
rect 12440 31977 12449 32011
rect 12449 31977 12483 32011
rect 12483 31977 12492 32011
rect 12440 31968 12492 31977
rect 12992 32011 13044 32020
rect 12992 31977 13001 32011
rect 13001 31977 13035 32011
rect 13035 31977 13044 32011
rect 12992 31968 13044 31977
rect 15200 31968 15252 32020
rect 20168 31968 20220 32020
rect 20260 31968 20312 32020
rect 21272 31968 21324 32020
rect 26516 31968 26568 32020
rect 26700 31968 26752 32020
rect 30472 32011 30524 32020
rect 30472 31977 30481 32011
rect 30481 31977 30515 32011
rect 30515 31977 30524 32011
rect 30472 31968 30524 31977
rect 30748 31968 30800 32020
rect 3884 31900 3936 31952
rect 3148 31875 3200 31884
rect 3148 31841 3157 31875
rect 3157 31841 3191 31875
rect 3191 31841 3200 31875
rect 3148 31832 3200 31841
rect 4528 31875 4580 31884
rect 4528 31841 4537 31875
rect 4537 31841 4571 31875
rect 4571 31841 4580 31875
rect 4528 31832 4580 31841
rect 5724 31832 5776 31884
rect 6828 31900 6880 31952
rect 7288 31900 7340 31952
rect 11152 31900 11204 31952
rect 4344 31807 4396 31816
rect 4344 31773 4353 31807
rect 4353 31773 4387 31807
rect 4387 31773 4396 31807
rect 4344 31764 4396 31773
rect 5448 31807 5500 31816
rect 5448 31773 5457 31807
rect 5457 31773 5491 31807
rect 5491 31773 5500 31807
rect 5448 31764 5500 31773
rect 10416 31832 10468 31884
rect 14372 31900 14424 31952
rect 17408 31900 17460 31952
rect 21916 31900 21968 31952
rect 29276 31900 29328 31952
rect 30012 31900 30064 31952
rect 15108 31875 15160 31884
rect 9864 31764 9916 31816
rect 15108 31841 15117 31875
rect 15117 31841 15151 31875
rect 15151 31841 15160 31875
rect 15108 31832 15160 31841
rect 16304 31832 16356 31884
rect 23020 31832 23072 31884
rect 25872 31875 25924 31884
rect 25872 31841 25881 31875
rect 25881 31841 25915 31875
rect 25915 31841 25924 31875
rect 25872 31832 25924 31841
rect 29552 31832 29604 31884
rect 5724 31696 5776 31748
rect 9680 31696 9732 31748
rect 10048 31696 10100 31748
rect 7196 31628 7248 31680
rect 12808 31696 12860 31748
rect 13176 31696 13228 31748
rect 12532 31628 12584 31680
rect 16580 31807 16632 31816
rect 16580 31773 16589 31807
rect 16589 31773 16623 31807
rect 16623 31773 16632 31807
rect 16580 31764 16632 31773
rect 22100 31764 22152 31816
rect 23572 31764 23624 31816
rect 29460 31764 29512 31816
rect 29920 31764 29972 31816
rect 20720 31696 20772 31748
rect 29368 31696 29420 31748
rect 30656 31696 30708 31748
rect 17960 31628 18012 31680
rect 28080 31628 28132 31680
rect 31208 31764 31260 31816
rect 31668 31764 31720 31816
rect 6517 31526 6569 31578
rect 6581 31526 6633 31578
rect 6645 31526 6697 31578
rect 6709 31526 6761 31578
rect 17588 31526 17640 31578
rect 17652 31526 17704 31578
rect 17716 31526 17768 31578
rect 17780 31526 17832 31578
rect 28658 31526 28710 31578
rect 28722 31526 28774 31578
rect 28786 31526 28838 31578
rect 28850 31526 28902 31578
rect 3148 31288 3200 31340
rect 3700 31288 3752 31340
rect 4344 31356 4396 31408
rect 4988 31288 5040 31340
rect 5356 31288 5408 31340
rect 5540 31220 5592 31272
rect 7380 31220 7432 31272
rect 9956 31220 10008 31272
rect 15108 31424 15160 31476
rect 16580 31424 16632 31476
rect 20720 31424 20772 31476
rect 12532 31331 12584 31340
rect 12532 31297 12541 31331
rect 12541 31297 12575 31331
rect 12575 31297 12584 31331
rect 12532 31288 12584 31297
rect 9772 31152 9824 31204
rect 9864 31152 9916 31204
rect 11612 31220 11664 31272
rect 13360 31220 13412 31272
rect 13912 31263 13964 31272
rect 13912 31229 13921 31263
rect 13921 31229 13955 31263
rect 13955 31229 13964 31263
rect 13912 31220 13964 31229
rect 16120 31220 16172 31272
rect 15292 31152 15344 31204
rect 18144 31331 18196 31340
rect 18144 31297 18153 31331
rect 18153 31297 18187 31331
rect 18187 31297 18196 31331
rect 18144 31288 18196 31297
rect 18604 31288 18656 31340
rect 23572 31331 23624 31340
rect 17960 31263 18012 31272
rect 17960 31229 17969 31263
rect 17969 31229 18003 31263
rect 18003 31229 18012 31263
rect 23572 31297 23581 31331
rect 23581 31297 23615 31331
rect 23615 31297 23624 31331
rect 23572 31288 23624 31297
rect 24308 31288 24360 31340
rect 28080 31331 28132 31340
rect 22836 31263 22888 31272
rect 17960 31220 18012 31229
rect 22836 31229 22845 31263
rect 22845 31229 22879 31263
rect 22879 31229 22888 31263
rect 22836 31220 22888 31229
rect 23940 31263 23992 31272
rect 23940 31229 23949 31263
rect 23949 31229 23983 31263
rect 23983 31229 23992 31263
rect 23940 31220 23992 31229
rect 3148 31084 3200 31136
rect 5908 31084 5960 31136
rect 7104 31084 7156 31136
rect 8208 31084 8260 31136
rect 10140 31127 10192 31136
rect 10140 31093 10149 31127
rect 10149 31093 10183 31127
rect 10183 31093 10192 31127
rect 10140 31084 10192 31093
rect 12440 31084 12492 31136
rect 13084 31127 13136 31136
rect 13084 31093 13093 31127
rect 13093 31093 13127 31127
rect 13127 31093 13136 31127
rect 13084 31084 13136 31093
rect 14372 31127 14424 31136
rect 14372 31093 14381 31127
rect 14381 31093 14415 31127
rect 14415 31093 14424 31127
rect 14372 31084 14424 31093
rect 19616 31152 19668 31204
rect 28080 31297 28089 31331
rect 28089 31297 28123 31331
rect 28123 31297 28132 31331
rect 28080 31288 28132 31297
rect 31300 31288 31352 31340
rect 27620 31220 27672 31272
rect 27804 31263 27856 31272
rect 27804 31229 27813 31263
rect 27813 31229 27847 31263
rect 27847 31229 27856 31263
rect 27804 31220 27856 31229
rect 31668 31220 31720 31272
rect 26516 31152 26568 31204
rect 29368 31152 29420 31204
rect 17960 31084 18012 31136
rect 19064 31084 19116 31136
rect 25320 31084 25372 31136
rect 29552 31127 29604 31136
rect 29552 31093 29561 31127
rect 29561 31093 29595 31127
rect 29595 31093 29604 31127
rect 29552 31084 29604 31093
rect 31024 31084 31076 31136
rect 31300 31127 31352 31136
rect 31300 31093 31309 31127
rect 31309 31093 31343 31127
rect 31343 31093 31352 31127
rect 31300 31084 31352 31093
rect 12052 30982 12104 31034
rect 12116 30982 12168 31034
rect 12180 30982 12232 31034
rect 12244 30982 12296 31034
rect 23123 30982 23175 31034
rect 23187 30982 23239 31034
rect 23251 30982 23303 31034
rect 23315 30982 23367 31034
rect 6828 30880 6880 30932
rect 11612 30923 11664 30932
rect 11612 30889 11621 30923
rect 11621 30889 11655 30923
rect 11655 30889 11664 30923
rect 11612 30880 11664 30889
rect 12440 30923 12492 30932
rect 12440 30889 12449 30923
rect 12449 30889 12483 30923
rect 12483 30889 12492 30923
rect 12440 30880 12492 30889
rect 13912 30880 13964 30932
rect 14924 30880 14976 30932
rect 17960 30880 18012 30932
rect 23480 30880 23532 30932
rect 23940 30880 23992 30932
rect 25320 30880 25372 30932
rect 30656 30880 30708 30932
rect 5448 30812 5500 30864
rect 3148 30787 3200 30796
rect 3148 30753 3157 30787
rect 3157 30753 3191 30787
rect 3191 30753 3200 30787
rect 3148 30744 3200 30753
rect 4804 30744 4856 30796
rect 5632 30787 5684 30796
rect 5632 30753 5641 30787
rect 5641 30753 5675 30787
rect 5675 30753 5684 30787
rect 5632 30744 5684 30753
rect 5908 30787 5960 30796
rect 5908 30753 5917 30787
rect 5917 30753 5951 30787
rect 5951 30753 5960 30787
rect 5908 30744 5960 30753
rect 17408 30812 17460 30864
rect 31668 30880 31720 30932
rect 7104 30787 7156 30796
rect 7104 30753 7113 30787
rect 7113 30753 7147 30787
rect 7147 30753 7156 30787
rect 7104 30744 7156 30753
rect 10048 30744 10100 30796
rect 12624 30744 12676 30796
rect 13636 30744 13688 30796
rect 14372 30744 14424 30796
rect 20536 30787 20588 30796
rect 20536 30753 20545 30787
rect 20545 30753 20579 30787
rect 20579 30753 20588 30787
rect 20536 30744 20588 30753
rect 22836 30787 22888 30796
rect 22836 30753 22845 30787
rect 22845 30753 22879 30787
rect 22879 30753 22888 30787
rect 23940 30787 23992 30796
rect 22836 30744 22888 30753
rect 2964 30719 3016 30728
rect 2964 30685 2973 30719
rect 2973 30685 3007 30719
rect 3007 30685 3016 30719
rect 2964 30676 3016 30685
rect 3056 30719 3108 30728
rect 3056 30685 3065 30719
rect 3065 30685 3099 30719
rect 3099 30685 3108 30719
rect 3240 30719 3292 30728
rect 3056 30676 3108 30685
rect 3240 30685 3249 30719
rect 3249 30685 3283 30719
rect 3283 30685 3292 30719
rect 3240 30676 3292 30685
rect 4988 30719 5040 30728
rect 4988 30685 4997 30719
rect 4997 30685 5031 30719
rect 5031 30685 5040 30719
rect 4988 30676 5040 30685
rect 7012 30719 7064 30728
rect 2780 30583 2832 30592
rect 2780 30549 2789 30583
rect 2789 30549 2823 30583
rect 2823 30549 2832 30583
rect 4068 30608 4120 30660
rect 5724 30608 5776 30660
rect 7012 30685 7021 30719
rect 7021 30685 7055 30719
rect 7055 30685 7064 30719
rect 7012 30676 7064 30685
rect 9956 30676 10008 30728
rect 13360 30676 13412 30728
rect 16120 30719 16172 30728
rect 16120 30685 16129 30719
rect 16129 30685 16163 30719
rect 16163 30685 16172 30719
rect 16120 30676 16172 30685
rect 17408 30676 17460 30728
rect 19616 30676 19668 30728
rect 20352 30608 20404 30660
rect 23940 30753 23949 30787
rect 23949 30753 23983 30787
rect 23983 30753 23992 30787
rect 23940 30744 23992 30753
rect 26516 30812 26568 30864
rect 31024 30855 31076 30864
rect 31024 30821 31033 30855
rect 31033 30821 31067 30855
rect 31067 30821 31076 30855
rect 31024 30812 31076 30821
rect 31484 30812 31536 30864
rect 27620 30744 27672 30796
rect 26240 30676 26292 30728
rect 27344 30719 27396 30728
rect 27344 30685 27353 30719
rect 27353 30685 27387 30719
rect 27387 30685 27396 30719
rect 27344 30676 27396 30685
rect 24860 30608 24912 30660
rect 2780 30540 2832 30549
rect 10876 30540 10928 30592
rect 21088 30540 21140 30592
rect 6517 30438 6569 30490
rect 6581 30438 6633 30490
rect 6645 30438 6697 30490
rect 6709 30438 6761 30490
rect 17588 30438 17640 30490
rect 17652 30438 17704 30490
rect 17716 30438 17768 30490
rect 17780 30438 17832 30490
rect 28658 30438 28710 30490
rect 28722 30438 28774 30490
rect 28786 30438 28838 30490
rect 28850 30438 28902 30490
rect 4804 30379 4856 30388
rect 4804 30345 4813 30379
rect 4813 30345 4847 30379
rect 4847 30345 4856 30379
rect 10048 30379 10100 30388
rect 4804 30336 4856 30345
rect 10048 30345 10057 30379
rect 10057 30345 10091 30379
rect 10091 30345 10100 30379
rect 10048 30336 10100 30345
rect 7012 30268 7064 30320
rect 7472 30243 7524 30252
rect 7472 30209 7481 30243
rect 7481 30209 7515 30243
rect 7515 30209 7524 30243
rect 7472 30200 7524 30209
rect 1400 30175 1452 30184
rect 1400 30141 1409 30175
rect 1409 30141 1443 30175
rect 1443 30141 1452 30175
rect 1400 30132 1452 30141
rect 2780 30132 2832 30184
rect 3700 30175 3752 30184
rect 3700 30141 3709 30175
rect 3709 30141 3743 30175
rect 3743 30141 3752 30175
rect 3700 30132 3752 30141
rect 4252 30132 4304 30184
rect 8208 30132 8260 30184
rect 10140 30175 10192 30184
rect 5724 30064 5776 30116
rect 10140 30141 10149 30175
rect 10149 30141 10183 30175
rect 10183 30141 10192 30175
rect 10140 30132 10192 30141
rect 10600 30175 10652 30184
rect 10600 30141 10609 30175
rect 10609 30141 10643 30175
rect 10643 30141 10652 30175
rect 10600 30132 10652 30141
rect 10968 30132 11020 30184
rect 12440 30132 12492 30184
rect 12992 30132 13044 30184
rect 11612 30064 11664 30116
rect 15292 30268 15344 30320
rect 17408 30268 17460 30320
rect 17960 30200 18012 30252
rect 19156 30200 19208 30252
rect 20352 30200 20404 30252
rect 21088 30243 21140 30252
rect 21088 30209 21097 30243
rect 21097 30209 21131 30243
rect 21131 30209 21140 30243
rect 21088 30200 21140 30209
rect 23572 30336 23624 30388
rect 23940 30336 23992 30388
rect 24768 30336 24820 30388
rect 27344 30268 27396 30320
rect 14188 30175 14240 30184
rect 14188 30141 14197 30175
rect 14197 30141 14231 30175
rect 14231 30141 14240 30175
rect 14188 30132 14240 30141
rect 14924 30175 14976 30184
rect 14924 30141 14933 30175
rect 14933 30141 14967 30175
rect 14967 30141 14976 30175
rect 14924 30132 14976 30141
rect 18604 30175 18656 30184
rect 13912 30064 13964 30116
rect 3148 29996 3200 30048
rect 8576 29996 8628 30048
rect 10876 29996 10928 30048
rect 12808 29996 12860 30048
rect 12992 29996 13044 30048
rect 18604 30141 18613 30175
rect 18613 30141 18647 30175
rect 18647 30141 18656 30175
rect 18604 30132 18656 30141
rect 20996 30132 21048 30184
rect 21364 30132 21416 30184
rect 23480 30200 23532 30252
rect 26608 30243 26660 30252
rect 26608 30209 26617 30243
rect 26617 30209 26651 30243
rect 26651 30209 26660 30243
rect 26608 30200 26660 30209
rect 28356 30200 28408 30252
rect 24860 30132 24912 30184
rect 26148 30132 26200 30184
rect 26240 30132 26292 30184
rect 29552 30132 29604 30184
rect 29920 30200 29972 30252
rect 30012 30175 30064 30184
rect 30012 30141 30021 30175
rect 30021 30141 30055 30175
rect 30055 30141 30064 30175
rect 30012 30132 30064 30141
rect 19616 29996 19668 30048
rect 24308 30064 24360 30116
rect 21180 29996 21232 30048
rect 25872 29996 25924 30048
rect 26424 30039 26476 30048
rect 26424 30005 26433 30039
rect 26433 30005 26467 30039
rect 26467 30005 26476 30039
rect 26424 29996 26476 30005
rect 12052 29894 12104 29946
rect 12116 29894 12168 29946
rect 12180 29894 12232 29946
rect 12244 29894 12296 29946
rect 23123 29894 23175 29946
rect 23187 29894 23239 29946
rect 23251 29894 23303 29946
rect 23315 29894 23367 29946
rect 3240 29792 3292 29844
rect 5632 29835 5684 29844
rect 5632 29801 5641 29835
rect 5641 29801 5675 29835
rect 5675 29801 5684 29835
rect 5632 29792 5684 29801
rect 9772 29835 9824 29844
rect 9772 29801 9781 29835
rect 9781 29801 9815 29835
rect 9815 29801 9824 29835
rect 9772 29792 9824 29801
rect 10968 29835 11020 29844
rect 10968 29801 10977 29835
rect 10977 29801 11011 29835
rect 11011 29801 11020 29835
rect 10968 29792 11020 29801
rect 13084 29792 13136 29844
rect 16120 29792 16172 29844
rect 3148 29699 3200 29708
rect 3148 29665 3157 29699
rect 3157 29665 3191 29699
rect 3191 29665 3200 29699
rect 3148 29656 3200 29665
rect 5724 29699 5776 29708
rect 5724 29665 5733 29699
rect 5733 29665 5767 29699
rect 5767 29665 5776 29699
rect 5724 29656 5776 29665
rect 5908 29699 5960 29708
rect 5908 29665 5917 29699
rect 5917 29665 5951 29699
rect 5951 29665 5960 29699
rect 5908 29656 5960 29665
rect 8024 29656 8076 29708
rect 8576 29656 8628 29708
rect 10232 29699 10284 29708
rect 10232 29665 10241 29699
rect 10241 29665 10275 29699
rect 10275 29665 10284 29699
rect 10232 29656 10284 29665
rect 4344 29588 4396 29640
rect 4988 29588 5040 29640
rect 7656 29631 7708 29640
rect 7656 29597 7665 29631
rect 7665 29597 7699 29631
rect 7699 29597 7708 29631
rect 7656 29588 7708 29597
rect 3424 29452 3476 29504
rect 9128 29452 9180 29504
rect 9864 29520 9916 29572
rect 10600 29656 10652 29708
rect 11428 29724 11480 29776
rect 12716 29724 12768 29776
rect 16396 29767 16448 29776
rect 16396 29733 16414 29767
rect 16414 29733 16448 29767
rect 16396 29724 16448 29733
rect 16764 29724 16816 29776
rect 11612 29631 11664 29640
rect 11612 29597 11621 29631
rect 11621 29597 11655 29631
rect 11655 29597 11664 29631
rect 11612 29588 11664 29597
rect 14372 29656 14424 29708
rect 12900 29588 12952 29640
rect 12440 29520 12492 29572
rect 16120 29656 16172 29708
rect 18420 29656 18472 29708
rect 21180 29792 21232 29844
rect 31760 29792 31812 29844
rect 24768 29656 24820 29708
rect 25504 29656 25556 29708
rect 26424 29724 26476 29776
rect 26240 29699 26292 29708
rect 26240 29665 26249 29699
rect 26249 29665 26283 29699
rect 26283 29665 26292 29699
rect 26240 29656 26292 29665
rect 17224 29631 17276 29640
rect 17224 29597 17233 29631
rect 17233 29597 17267 29631
rect 17267 29597 17276 29631
rect 17224 29588 17276 29597
rect 18328 29588 18380 29640
rect 18604 29588 18656 29640
rect 20904 29588 20956 29640
rect 21456 29631 21508 29640
rect 21456 29597 21465 29631
rect 21465 29597 21499 29631
rect 21499 29597 21508 29631
rect 21456 29588 21508 29597
rect 24860 29520 24912 29572
rect 26240 29520 26292 29572
rect 28356 29699 28408 29708
rect 28356 29665 28365 29699
rect 28365 29665 28399 29699
rect 28399 29665 28408 29699
rect 28356 29656 28408 29665
rect 29000 29656 29052 29708
rect 27620 29588 27672 29640
rect 30932 29631 30984 29640
rect 30932 29597 30941 29631
rect 30941 29597 30975 29631
rect 30975 29597 30984 29631
rect 30932 29588 30984 29597
rect 27896 29563 27948 29572
rect 27896 29529 27905 29563
rect 27905 29529 27939 29563
rect 27939 29529 27948 29563
rect 27896 29520 27948 29529
rect 12900 29452 12952 29504
rect 13728 29452 13780 29504
rect 16672 29452 16724 29504
rect 20536 29452 20588 29504
rect 22008 29452 22060 29504
rect 25136 29452 25188 29504
rect 31300 29452 31352 29504
rect 6517 29350 6569 29402
rect 6581 29350 6633 29402
rect 6645 29350 6697 29402
rect 6709 29350 6761 29402
rect 17588 29350 17640 29402
rect 17652 29350 17704 29402
rect 17716 29350 17768 29402
rect 17780 29350 17832 29402
rect 28658 29350 28710 29402
rect 28722 29350 28774 29402
rect 28786 29350 28838 29402
rect 28850 29350 28902 29402
rect 8024 29291 8076 29300
rect 4068 29180 4120 29232
rect 5448 29180 5500 29232
rect 3240 29155 3292 29164
rect 3240 29121 3249 29155
rect 3249 29121 3283 29155
rect 3283 29121 3292 29155
rect 3240 29112 3292 29121
rect 3424 29155 3476 29164
rect 3424 29121 3433 29155
rect 3433 29121 3467 29155
rect 3467 29121 3476 29155
rect 3424 29112 3476 29121
rect 7196 29112 7248 29164
rect 8024 29257 8033 29291
rect 8033 29257 8067 29291
rect 8067 29257 8076 29291
rect 8024 29248 8076 29257
rect 9864 29291 9916 29300
rect 9864 29257 9873 29291
rect 9873 29257 9907 29291
rect 9907 29257 9916 29291
rect 9864 29248 9916 29257
rect 12440 29291 12492 29300
rect 12440 29257 12449 29291
rect 12449 29257 12483 29291
rect 12483 29257 12492 29291
rect 12716 29291 12768 29300
rect 12440 29248 12492 29257
rect 12716 29257 12725 29291
rect 12725 29257 12759 29291
rect 12759 29257 12768 29291
rect 12716 29248 12768 29257
rect 18328 29291 18380 29300
rect 18328 29257 18337 29291
rect 18337 29257 18371 29291
rect 18371 29257 18380 29291
rect 18328 29248 18380 29257
rect 20904 29248 20956 29300
rect 25320 29291 25372 29300
rect 25320 29257 25329 29291
rect 25329 29257 25363 29291
rect 25363 29257 25372 29291
rect 25320 29248 25372 29257
rect 25504 29291 25556 29300
rect 25504 29257 25513 29291
rect 25513 29257 25547 29291
rect 25547 29257 25556 29291
rect 25504 29248 25556 29257
rect 30932 29248 30984 29300
rect 7656 29180 7708 29232
rect 8208 29112 8260 29164
rect 11888 29180 11940 29232
rect 12532 29180 12584 29232
rect 13176 29112 13228 29164
rect 27620 29180 27672 29232
rect 16672 29112 16724 29164
rect 1768 29087 1820 29096
rect 1768 29053 1777 29087
rect 1777 29053 1811 29087
rect 1811 29053 1820 29087
rect 1768 29044 1820 29053
rect 3056 29044 3108 29096
rect 3332 29087 3384 29096
rect 3332 29053 3341 29087
rect 3341 29053 3375 29087
rect 3375 29053 3384 29087
rect 3332 29044 3384 29053
rect 4252 29087 4304 29096
rect 4252 29053 4261 29087
rect 4261 29053 4295 29087
rect 4295 29053 4304 29087
rect 4252 29044 4304 29053
rect 4344 29087 4396 29096
rect 4344 29053 4353 29087
rect 4353 29053 4387 29087
rect 4387 29053 4396 29087
rect 4344 29044 4396 29053
rect 3056 28951 3108 28960
rect 3056 28917 3065 28951
rect 3065 28917 3099 28951
rect 3099 28917 3108 28951
rect 3056 28908 3108 28917
rect 5080 28951 5132 28960
rect 5080 28917 5089 28951
rect 5089 28917 5123 28951
rect 5123 28917 5132 28951
rect 5080 28908 5132 28917
rect 5724 29044 5776 29096
rect 7656 29087 7708 29096
rect 7656 29053 7665 29087
rect 7665 29053 7699 29087
rect 7699 29053 7708 29087
rect 7656 29044 7708 29053
rect 9496 29044 9548 29096
rect 9956 29044 10008 29096
rect 10692 29087 10744 29096
rect 10692 29053 10701 29087
rect 10701 29053 10735 29087
rect 10735 29053 10744 29087
rect 10692 29044 10744 29053
rect 12900 29044 12952 29096
rect 13084 29087 13136 29096
rect 13084 29053 13093 29087
rect 13093 29053 13127 29087
rect 13127 29053 13136 29087
rect 13084 29044 13136 29053
rect 16764 29044 16816 29096
rect 18604 29112 18656 29164
rect 19156 29112 19208 29164
rect 19616 29044 19668 29096
rect 20444 29044 20496 29096
rect 20536 29087 20588 29096
rect 20536 29053 20545 29087
rect 20545 29053 20579 29087
rect 20579 29053 20588 29087
rect 24584 29112 24636 29164
rect 32404 29180 32456 29232
rect 31208 29155 31260 29164
rect 31208 29121 31217 29155
rect 31217 29121 31251 29155
rect 31251 29121 31260 29155
rect 31208 29112 31260 29121
rect 20536 29044 20588 29053
rect 5540 28976 5592 29028
rect 6828 28976 6880 29028
rect 12716 28976 12768 29028
rect 17408 28976 17460 29028
rect 22560 28976 22612 29028
rect 29368 29044 29420 29096
rect 30104 29044 30156 29096
rect 31300 29044 31352 29096
rect 33600 29087 33652 29096
rect 33600 29053 33609 29087
rect 33609 29053 33643 29087
rect 33643 29053 33652 29087
rect 33600 29044 33652 29053
rect 25136 29019 25188 29028
rect 25136 28985 25145 29019
rect 25145 28985 25179 29019
rect 25179 28985 25188 29019
rect 25136 28976 25188 28985
rect 28264 29019 28316 29028
rect 28264 28985 28273 29019
rect 28273 28985 28307 29019
rect 28307 28985 28316 29019
rect 28264 28976 28316 28985
rect 8852 28951 8904 28960
rect 8852 28917 8861 28951
rect 8861 28917 8895 28951
rect 8895 28917 8904 28951
rect 8852 28908 8904 28917
rect 10968 28908 11020 28960
rect 14556 28951 14608 28960
rect 14556 28917 14565 28951
rect 14565 28917 14599 28951
rect 14599 28917 14608 28951
rect 14556 28908 14608 28917
rect 14648 28951 14700 28960
rect 14648 28917 14657 28951
rect 14657 28917 14691 28951
rect 14691 28917 14700 28951
rect 15016 28951 15068 28960
rect 14648 28908 14700 28917
rect 15016 28917 15025 28951
rect 15025 28917 15059 28951
rect 15059 28917 15068 28951
rect 15016 28908 15068 28917
rect 20352 28951 20404 28960
rect 20352 28917 20361 28951
rect 20361 28917 20395 28951
rect 20395 28917 20404 28951
rect 20352 28908 20404 28917
rect 24308 28951 24360 28960
rect 24308 28917 24317 28951
rect 24317 28917 24351 28951
rect 24351 28917 24360 28951
rect 24308 28908 24360 28917
rect 25596 28908 25648 28960
rect 30288 28976 30340 29028
rect 12052 28806 12104 28858
rect 12116 28806 12168 28858
rect 12180 28806 12232 28858
rect 12244 28806 12296 28858
rect 23123 28806 23175 28858
rect 23187 28806 23239 28858
rect 23251 28806 23303 28858
rect 23315 28806 23367 28858
rect 4252 28704 4304 28756
rect 5724 28704 5776 28756
rect 8852 28704 8904 28756
rect 9128 28704 9180 28756
rect 10232 28747 10284 28756
rect 10232 28713 10241 28747
rect 10241 28713 10275 28747
rect 10275 28713 10284 28747
rect 10232 28704 10284 28713
rect 3056 28636 3108 28688
rect 5080 28679 5132 28688
rect 5080 28645 5114 28679
rect 5114 28645 5132 28679
rect 5080 28636 5132 28645
rect 10692 28636 10744 28688
rect 14556 28704 14608 28756
rect 14648 28704 14700 28756
rect 19340 28636 19392 28688
rect 21456 28704 21508 28756
rect 23480 28704 23532 28756
rect 25320 28704 25372 28756
rect 26332 28704 26384 28756
rect 28264 28704 28316 28756
rect 29000 28704 29052 28756
rect 1400 28568 1452 28620
rect 3884 28568 3936 28620
rect 8300 28568 8352 28620
rect 8576 28611 8628 28620
rect 5908 28500 5960 28552
rect 7472 28500 7524 28552
rect 8576 28577 8585 28611
rect 8585 28577 8619 28611
rect 8619 28577 8628 28611
rect 8576 28568 8628 28577
rect 9680 28568 9732 28620
rect 9864 28611 9916 28620
rect 9864 28577 9873 28611
rect 9873 28577 9907 28611
rect 9907 28577 9916 28611
rect 9864 28568 9916 28577
rect 10876 28568 10928 28620
rect 11060 28568 11112 28620
rect 12808 28611 12860 28620
rect 12808 28577 12817 28611
rect 12817 28577 12851 28611
rect 12851 28577 12860 28611
rect 12808 28568 12860 28577
rect 12992 28611 13044 28620
rect 12992 28577 13001 28611
rect 13001 28577 13035 28611
rect 13035 28577 13044 28611
rect 12992 28568 13044 28577
rect 13636 28611 13688 28620
rect 13636 28577 13645 28611
rect 13645 28577 13679 28611
rect 13679 28577 13688 28611
rect 13636 28568 13688 28577
rect 14004 28568 14056 28620
rect 16764 28611 16816 28620
rect 16764 28577 16773 28611
rect 16773 28577 16807 28611
rect 16807 28577 16816 28611
rect 16764 28568 16816 28577
rect 19064 28611 19116 28620
rect 19064 28577 19073 28611
rect 19073 28577 19107 28611
rect 19107 28577 19116 28611
rect 19064 28568 19116 28577
rect 20260 28611 20312 28620
rect 20260 28577 20269 28611
rect 20269 28577 20303 28611
rect 20303 28577 20312 28611
rect 20260 28568 20312 28577
rect 10048 28500 10100 28552
rect 13360 28432 13412 28484
rect 16672 28500 16724 28552
rect 20352 28500 20404 28552
rect 18972 28475 19024 28484
rect 18972 28441 18981 28475
rect 18981 28441 19015 28475
rect 19015 28441 19024 28475
rect 18972 28432 19024 28441
rect 20996 28611 21048 28620
rect 20996 28577 21005 28611
rect 21005 28577 21039 28611
rect 21039 28577 21048 28611
rect 20996 28568 21048 28577
rect 22008 28611 22060 28620
rect 22008 28577 22017 28611
rect 22017 28577 22051 28611
rect 22051 28577 22060 28611
rect 22008 28568 22060 28577
rect 22560 28568 22612 28620
rect 24768 28636 24820 28688
rect 26516 28636 26568 28688
rect 30288 28636 30340 28688
rect 32404 28679 32456 28688
rect 32404 28645 32438 28679
rect 32438 28645 32456 28679
rect 32404 28636 32456 28645
rect 24308 28568 24360 28620
rect 27620 28568 27672 28620
rect 21088 28543 21140 28552
rect 21088 28509 21097 28543
rect 21097 28509 21131 28543
rect 21131 28509 21140 28543
rect 21088 28500 21140 28509
rect 23940 28432 23992 28484
rect 6276 28364 6328 28416
rect 12624 28364 12676 28416
rect 16948 28407 17000 28416
rect 16948 28373 16957 28407
rect 16957 28373 16991 28407
rect 16991 28373 17000 28407
rect 16948 28364 17000 28373
rect 19340 28364 19392 28416
rect 22836 28364 22888 28416
rect 25780 28500 25832 28552
rect 29276 28543 29328 28552
rect 29276 28509 29285 28543
rect 29285 28509 29319 28543
rect 29319 28509 29328 28543
rect 29276 28500 29328 28509
rect 30288 28500 30340 28552
rect 31300 28500 31352 28552
rect 31944 28500 31996 28552
rect 31208 28432 31260 28484
rect 24124 28364 24176 28416
rect 25228 28364 25280 28416
rect 25688 28364 25740 28416
rect 33508 28407 33560 28416
rect 33508 28373 33517 28407
rect 33517 28373 33551 28407
rect 33551 28373 33560 28407
rect 33508 28364 33560 28373
rect 6517 28262 6569 28314
rect 6581 28262 6633 28314
rect 6645 28262 6697 28314
rect 6709 28262 6761 28314
rect 17588 28262 17640 28314
rect 17652 28262 17704 28314
rect 17716 28262 17768 28314
rect 17780 28262 17832 28314
rect 28658 28262 28710 28314
rect 28722 28262 28774 28314
rect 28786 28262 28838 28314
rect 28850 28262 28902 28314
rect 3332 28160 3384 28212
rect 4436 28203 4488 28212
rect 4436 28169 4445 28203
rect 4445 28169 4479 28203
rect 4479 28169 4488 28203
rect 4436 28160 4488 28169
rect 5540 28203 5592 28212
rect 5540 28169 5549 28203
rect 5549 28169 5583 28203
rect 5583 28169 5592 28203
rect 5540 28160 5592 28169
rect 11060 28203 11112 28212
rect 11060 28169 11069 28203
rect 11069 28169 11103 28203
rect 11103 28169 11112 28203
rect 11060 28160 11112 28169
rect 13912 28160 13964 28212
rect 21088 28160 21140 28212
rect 25780 28203 25832 28212
rect 25780 28169 25789 28203
rect 25789 28169 25823 28203
rect 25823 28169 25832 28203
rect 25780 28160 25832 28169
rect 29276 28160 29328 28212
rect 17316 28092 17368 28144
rect 9496 28024 9548 28076
rect 13728 28024 13780 28076
rect 16948 28024 17000 28076
rect 19156 28067 19208 28076
rect 19156 28033 19165 28067
rect 19165 28033 19199 28067
rect 19199 28033 19208 28067
rect 19156 28024 19208 28033
rect 25688 28135 25740 28144
rect 25688 28101 25697 28135
rect 25697 28101 25731 28135
rect 25731 28101 25740 28135
rect 25688 28092 25740 28101
rect 6276 27956 6328 28008
rect 8208 27956 8260 28008
rect 8392 27956 8444 28008
rect 10232 27999 10284 28008
rect 2964 27888 3016 27940
rect 4344 27931 4396 27940
rect 4344 27897 4353 27931
rect 4353 27897 4387 27931
rect 4387 27897 4396 27931
rect 4344 27888 4396 27897
rect 10232 27965 10241 27999
rect 10241 27965 10275 27999
rect 10275 27965 10284 27999
rect 10232 27956 10284 27965
rect 10968 27999 11020 28008
rect 10968 27965 10977 27999
rect 10977 27965 11011 27999
rect 11011 27965 11020 27999
rect 10968 27956 11020 27965
rect 12624 27956 12676 28008
rect 10140 27888 10192 27940
rect 12348 27888 12400 27940
rect 13084 27956 13136 28008
rect 15016 27956 15068 28008
rect 20260 28024 20312 28076
rect 20444 28024 20496 28076
rect 20812 27999 20864 28008
rect 20812 27965 20821 27999
rect 20821 27965 20855 27999
rect 20855 27965 20864 27999
rect 20812 27956 20864 27965
rect 21088 27956 21140 28008
rect 24860 28024 24912 28076
rect 17960 27931 18012 27940
rect 17960 27897 17969 27931
rect 17969 27897 18003 27931
rect 18003 27897 18012 27931
rect 17960 27888 18012 27897
rect 20720 27888 20772 27940
rect 8208 27863 8260 27872
rect 8208 27829 8217 27863
rect 8217 27829 8251 27863
rect 8251 27829 8260 27863
rect 8208 27820 8260 27829
rect 14188 27863 14240 27872
rect 14188 27829 14197 27863
rect 14197 27829 14231 27863
rect 14231 27829 14240 27863
rect 14188 27820 14240 27829
rect 14556 27863 14608 27872
rect 14556 27829 14565 27863
rect 14565 27829 14599 27863
rect 14599 27829 14608 27863
rect 14556 27820 14608 27829
rect 17408 27820 17460 27872
rect 18512 27863 18564 27872
rect 18512 27829 18521 27863
rect 18521 27829 18555 27863
rect 18555 27829 18564 27863
rect 18512 27820 18564 27829
rect 19064 27820 19116 27872
rect 19156 27820 19208 27872
rect 21180 27820 21232 27872
rect 22560 27888 22612 27940
rect 22836 27820 22888 27872
rect 23572 27820 23624 27872
rect 24032 27956 24084 28008
rect 24768 27999 24820 28008
rect 24768 27965 24777 27999
rect 24777 27965 24811 27999
rect 24811 27965 24820 27999
rect 24768 27956 24820 27965
rect 25320 27956 25372 28008
rect 27620 28024 27672 28076
rect 26332 27999 26384 28008
rect 26332 27965 26341 27999
rect 26341 27965 26375 27999
rect 26375 27965 26384 27999
rect 26332 27956 26384 27965
rect 26608 27956 26660 28008
rect 31208 28160 31260 28212
rect 26056 27888 26108 27940
rect 28724 27931 28776 27940
rect 28724 27897 28733 27931
rect 28733 27897 28767 27931
rect 28767 27897 28776 27931
rect 28724 27888 28776 27897
rect 30104 27888 30156 27940
rect 30380 27888 30432 27940
rect 25780 27820 25832 27872
rect 30656 27863 30708 27872
rect 30656 27829 30665 27863
rect 30665 27829 30699 27863
rect 30699 27829 30708 27863
rect 30656 27820 30708 27829
rect 12052 27718 12104 27770
rect 12116 27718 12168 27770
rect 12180 27718 12232 27770
rect 12244 27718 12296 27770
rect 23123 27718 23175 27770
rect 23187 27718 23239 27770
rect 23251 27718 23303 27770
rect 23315 27718 23367 27770
rect 4252 27616 4304 27668
rect 12992 27616 13044 27668
rect 14556 27616 14608 27668
rect 15016 27616 15068 27668
rect 20996 27659 21048 27668
rect 20996 27625 21005 27659
rect 21005 27625 21039 27659
rect 21039 27625 21048 27659
rect 20996 27616 21048 27625
rect 10140 27548 10192 27600
rect 10416 27591 10468 27600
rect 10416 27557 10425 27591
rect 10425 27557 10459 27591
rect 10459 27557 10468 27591
rect 10416 27548 10468 27557
rect 11428 27591 11480 27600
rect 11428 27557 11437 27591
rect 11437 27557 11471 27591
rect 11471 27557 11480 27591
rect 11428 27548 11480 27557
rect 14188 27548 14240 27600
rect 18420 27548 18472 27600
rect 20720 27591 20772 27600
rect 20720 27557 20729 27591
rect 20729 27557 20763 27591
rect 20763 27557 20772 27591
rect 20720 27548 20772 27557
rect 22100 27616 22152 27668
rect 25228 27659 25280 27668
rect 25228 27625 25237 27659
rect 25237 27625 25271 27659
rect 25271 27625 25280 27659
rect 25228 27616 25280 27625
rect 28724 27616 28776 27668
rect 33508 27616 33560 27668
rect 2964 27523 3016 27532
rect 2964 27489 2973 27523
rect 2973 27489 3007 27523
rect 3007 27489 3016 27523
rect 2964 27480 3016 27489
rect 2780 27412 2832 27464
rect 3148 27455 3200 27464
rect 3148 27421 3157 27455
rect 3157 27421 3191 27455
rect 3191 27421 3200 27455
rect 3148 27412 3200 27421
rect 4988 27412 5040 27464
rect 6092 27387 6144 27396
rect 6092 27353 6101 27387
rect 6101 27353 6135 27387
rect 6135 27353 6144 27387
rect 6092 27344 6144 27353
rect 2688 27319 2740 27328
rect 2688 27285 2697 27319
rect 2697 27285 2731 27319
rect 2731 27285 2740 27319
rect 2688 27276 2740 27285
rect 4528 27276 4580 27328
rect 7288 27276 7340 27328
rect 8392 27523 8444 27532
rect 8392 27489 8401 27523
rect 8401 27489 8435 27523
rect 8435 27489 8444 27523
rect 8392 27480 8444 27489
rect 9956 27480 10008 27532
rect 10232 27523 10284 27532
rect 10232 27489 10241 27523
rect 10241 27489 10275 27523
rect 10275 27489 10284 27523
rect 10232 27480 10284 27489
rect 11244 27480 11296 27532
rect 11520 27523 11572 27532
rect 11520 27489 11529 27523
rect 11529 27489 11563 27523
rect 11563 27489 11572 27523
rect 11520 27480 11572 27489
rect 11704 27480 11756 27532
rect 12440 27480 12492 27532
rect 13452 27523 13504 27532
rect 13452 27489 13461 27523
rect 13461 27489 13495 27523
rect 13495 27489 13504 27523
rect 13452 27480 13504 27489
rect 15016 27480 15068 27532
rect 17224 27523 17276 27532
rect 8760 27412 8812 27464
rect 10048 27412 10100 27464
rect 11060 27412 11112 27464
rect 11612 27412 11664 27464
rect 14740 27412 14792 27464
rect 17224 27489 17233 27523
rect 17233 27489 17267 27523
rect 17267 27489 17276 27523
rect 17224 27480 17276 27489
rect 19432 27480 19484 27532
rect 19800 27480 19852 27532
rect 20812 27480 20864 27532
rect 18512 27412 18564 27464
rect 21088 27480 21140 27532
rect 33324 27548 33376 27600
rect 22376 27523 22428 27532
rect 22376 27489 22385 27523
rect 22385 27489 22419 27523
rect 22419 27489 22428 27523
rect 22376 27480 22428 27489
rect 22468 27523 22520 27532
rect 22468 27489 22477 27523
rect 22477 27489 22511 27523
rect 22511 27489 22520 27523
rect 22468 27480 22520 27489
rect 22100 27412 22152 27464
rect 25044 27480 25096 27532
rect 25136 27480 25188 27532
rect 26240 27480 26292 27532
rect 26700 27480 26752 27532
rect 28264 27480 28316 27532
rect 30656 27480 30708 27532
rect 31944 27455 31996 27464
rect 31944 27421 31953 27455
rect 31953 27421 31987 27455
rect 31987 27421 31996 27455
rect 31944 27412 31996 27421
rect 15108 27344 15160 27396
rect 24032 27344 24084 27396
rect 24584 27387 24636 27396
rect 24584 27353 24593 27387
rect 24593 27353 24627 27387
rect 24627 27353 24636 27387
rect 24584 27344 24636 27353
rect 26332 27344 26384 27396
rect 30472 27344 30524 27396
rect 12072 27319 12124 27328
rect 12072 27285 12081 27319
rect 12081 27285 12115 27319
rect 12115 27285 12124 27319
rect 12072 27276 12124 27285
rect 12348 27276 12400 27328
rect 19064 27276 19116 27328
rect 20168 27319 20220 27328
rect 20168 27285 20177 27319
rect 20177 27285 20211 27319
rect 20211 27285 20220 27319
rect 20168 27276 20220 27285
rect 22652 27276 22704 27328
rect 22744 27276 22796 27328
rect 30564 27319 30616 27328
rect 30564 27285 30573 27319
rect 30573 27285 30607 27319
rect 30607 27285 30616 27319
rect 30564 27276 30616 27285
rect 31208 27276 31260 27328
rect 32588 27319 32640 27328
rect 32588 27285 32597 27319
rect 32597 27285 32631 27319
rect 32631 27285 32640 27319
rect 32588 27276 32640 27285
rect 6517 27174 6569 27226
rect 6581 27174 6633 27226
rect 6645 27174 6697 27226
rect 6709 27174 6761 27226
rect 17588 27174 17640 27226
rect 17652 27174 17704 27226
rect 17716 27174 17768 27226
rect 17780 27174 17832 27226
rect 28658 27174 28710 27226
rect 28722 27174 28774 27226
rect 28786 27174 28838 27226
rect 28850 27174 28902 27226
rect 9864 27072 9916 27124
rect 11520 27072 11572 27124
rect 12348 27115 12400 27124
rect 12348 27081 12357 27115
rect 12357 27081 12391 27115
rect 12391 27081 12400 27115
rect 12348 27072 12400 27081
rect 13452 27115 13504 27124
rect 13452 27081 13461 27115
rect 13461 27081 13495 27115
rect 13495 27081 13504 27115
rect 13452 27072 13504 27081
rect 13544 27072 13596 27124
rect 11244 27004 11296 27056
rect 13084 27004 13136 27056
rect 1492 26979 1544 26988
rect 1492 26945 1501 26979
rect 1501 26945 1535 26979
rect 1535 26945 1544 26979
rect 1492 26936 1544 26945
rect 2688 26868 2740 26920
rect 4528 26911 4580 26920
rect 4528 26877 4537 26911
rect 4537 26877 4571 26911
rect 4571 26877 4580 26911
rect 4528 26868 4580 26877
rect 6092 26936 6144 26988
rect 7932 26979 7984 26988
rect 7932 26945 7941 26979
rect 7941 26945 7975 26979
rect 7975 26945 7984 26979
rect 7932 26936 7984 26945
rect 9036 26936 9088 26988
rect 13452 26936 13504 26988
rect 14188 26936 14240 26988
rect 8208 26868 8260 26920
rect 8668 26911 8720 26920
rect 8668 26877 8677 26911
rect 8677 26877 8711 26911
rect 8711 26877 8720 26911
rect 8668 26868 8720 26877
rect 8944 26911 8996 26920
rect 8944 26877 8953 26911
rect 8953 26877 8987 26911
rect 8987 26877 8996 26911
rect 8944 26868 8996 26877
rect 9496 26911 9548 26920
rect 9496 26877 9505 26911
rect 9505 26877 9539 26911
rect 9539 26877 9548 26911
rect 9496 26868 9548 26877
rect 10600 26911 10652 26920
rect 10600 26877 10609 26911
rect 10609 26877 10643 26911
rect 10643 26877 10652 26911
rect 10600 26868 10652 26877
rect 11152 26868 11204 26920
rect 12440 26911 12492 26920
rect 12440 26877 12449 26911
rect 12449 26877 12483 26911
rect 12483 26877 12492 26911
rect 12900 26911 12952 26920
rect 12440 26868 12492 26877
rect 12900 26877 12909 26911
rect 12909 26877 12943 26911
rect 12943 26877 12952 26911
rect 12900 26868 12952 26877
rect 13268 26911 13320 26920
rect 13268 26877 13277 26911
rect 13277 26877 13311 26911
rect 13311 26877 13320 26911
rect 13268 26868 13320 26877
rect 13820 26868 13872 26920
rect 20168 27072 20220 27124
rect 22192 27072 22244 27124
rect 22836 27072 22888 27124
rect 24768 27115 24820 27124
rect 22928 27004 22980 27056
rect 16672 26936 16724 26988
rect 17960 26936 18012 26988
rect 19432 26979 19484 26988
rect 19432 26945 19441 26979
rect 19441 26945 19475 26979
rect 19475 26945 19484 26979
rect 19432 26936 19484 26945
rect 20720 26936 20772 26988
rect 21180 26936 21232 26988
rect 22744 26979 22796 26988
rect 22744 26945 22753 26979
rect 22753 26945 22787 26979
rect 22787 26945 22796 26979
rect 22744 26936 22796 26945
rect 14924 26868 14976 26920
rect 16580 26868 16632 26920
rect 17316 26911 17368 26920
rect 17316 26877 17325 26911
rect 17325 26877 17359 26911
rect 17359 26877 17368 26911
rect 17316 26868 17368 26877
rect 4896 26800 4948 26852
rect 4988 26800 5040 26852
rect 2872 26775 2924 26784
rect 2872 26741 2881 26775
rect 2881 26741 2915 26775
rect 2915 26741 2924 26775
rect 2872 26732 2924 26741
rect 3332 26775 3384 26784
rect 3332 26741 3341 26775
rect 3341 26741 3375 26775
rect 3375 26741 3384 26775
rect 3332 26732 3384 26741
rect 10324 26800 10376 26852
rect 12072 26800 12124 26852
rect 18604 26868 18656 26920
rect 19064 26868 19116 26920
rect 22192 26868 22244 26920
rect 22652 26911 22704 26920
rect 22652 26877 22661 26911
rect 22661 26877 22695 26911
rect 22695 26877 22704 26911
rect 22652 26868 22704 26877
rect 23020 26868 23072 26920
rect 24768 27081 24777 27115
rect 24777 27081 24811 27115
rect 24811 27081 24820 27115
rect 24768 27072 24820 27081
rect 25044 27004 25096 27056
rect 27620 27004 27672 27056
rect 31760 27072 31812 27124
rect 25320 26936 25372 26988
rect 29828 26979 29880 26988
rect 29828 26945 29837 26979
rect 29837 26945 29871 26979
rect 29871 26945 29880 26979
rect 29828 26936 29880 26945
rect 24032 26911 24084 26920
rect 24032 26877 24041 26911
rect 24041 26877 24075 26911
rect 24075 26877 24084 26911
rect 24032 26868 24084 26877
rect 5908 26775 5960 26784
rect 5908 26741 5917 26775
rect 5917 26741 5951 26775
rect 5951 26741 5960 26775
rect 5908 26732 5960 26741
rect 7472 26775 7524 26784
rect 7472 26741 7481 26775
rect 7481 26741 7515 26775
rect 7515 26741 7524 26775
rect 7472 26732 7524 26741
rect 8760 26775 8812 26784
rect 8760 26741 8769 26775
rect 8769 26741 8803 26775
rect 8803 26741 8812 26775
rect 8760 26732 8812 26741
rect 13636 26732 13688 26784
rect 20444 26775 20496 26784
rect 20444 26741 20453 26775
rect 20453 26741 20487 26775
rect 20487 26741 20496 26775
rect 20444 26732 20496 26741
rect 21088 26732 21140 26784
rect 26240 26868 26292 26920
rect 27804 26868 27856 26920
rect 30104 26911 30156 26920
rect 30104 26877 30113 26911
rect 30113 26877 30147 26911
rect 30147 26877 30156 26911
rect 30104 26868 30156 26877
rect 33232 26936 33284 26988
rect 24860 26800 24912 26852
rect 31576 26800 31628 26852
rect 24952 26732 25004 26784
rect 28172 26732 28224 26784
rect 32956 26732 33008 26784
rect 12052 26630 12104 26682
rect 12116 26630 12168 26682
rect 12180 26630 12232 26682
rect 12244 26630 12296 26682
rect 23123 26630 23175 26682
rect 23187 26630 23239 26682
rect 23251 26630 23303 26682
rect 23315 26630 23367 26682
rect 3148 26528 3200 26580
rect 4896 26571 4948 26580
rect 4896 26537 4905 26571
rect 4905 26537 4939 26571
rect 4939 26537 4948 26571
rect 4896 26528 4948 26537
rect 7472 26571 7524 26580
rect 7472 26537 7481 26571
rect 7481 26537 7515 26571
rect 7515 26537 7524 26571
rect 7472 26528 7524 26537
rect 8392 26571 8444 26580
rect 8392 26537 8401 26571
rect 8401 26537 8435 26571
rect 8435 26537 8444 26571
rect 8392 26528 8444 26537
rect 10232 26528 10284 26580
rect 16580 26528 16632 26580
rect 18972 26528 19024 26580
rect 19432 26528 19484 26580
rect 20168 26528 20220 26580
rect 1584 26460 1636 26512
rect 10140 26460 10192 26512
rect 12164 26460 12216 26512
rect 12440 26503 12492 26512
rect 12440 26469 12470 26503
rect 12470 26469 12492 26503
rect 12440 26460 12492 26469
rect 13820 26460 13872 26512
rect 14740 26503 14792 26512
rect 14740 26469 14749 26503
rect 14749 26469 14783 26503
rect 14783 26469 14792 26503
rect 14740 26460 14792 26469
rect 16672 26503 16724 26512
rect 16672 26469 16681 26503
rect 16681 26469 16715 26503
rect 16715 26469 16724 26503
rect 16672 26460 16724 26469
rect 22928 26528 22980 26580
rect 25320 26528 25372 26580
rect 27804 26571 27856 26580
rect 27804 26537 27813 26571
rect 27813 26537 27847 26571
rect 27847 26537 27856 26571
rect 27804 26528 27856 26537
rect 33232 26528 33284 26580
rect 23020 26460 23072 26512
rect 26332 26503 26384 26512
rect 2872 26392 2924 26444
rect 4436 26392 4488 26444
rect 5080 26435 5132 26444
rect 5080 26401 5089 26435
rect 5089 26401 5123 26435
rect 5123 26401 5132 26435
rect 5080 26392 5132 26401
rect 5908 26392 5960 26444
rect 7932 26392 7984 26444
rect 10416 26435 10468 26444
rect 10416 26401 10425 26435
rect 10425 26401 10459 26435
rect 10459 26401 10468 26435
rect 10416 26392 10468 26401
rect 10600 26392 10652 26444
rect 4344 26324 4396 26376
rect 5540 26367 5592 26376
rect 5540 26333 5549 26367
rect 5549 26333 5583 26367
rect 5583 26333 5592 26367
rect 5540 26324 5592 26333
rect 7196 26367 7248 26376
rect 7196 26333 7205 26367
rect 7205 26333 7239 26367
rect 7239 26333 7248 26367
rect 7196 26324 7248 26333
rect 10876 26392 10928 26444
rect 11980 26392 12032 26444
rect 14556 26392 14608 26444
rect 15568 26435 15620 26444
rect 15568 26401 15577 26435
rect 15577 26401 15611 26435
rect 15611 26401 15620 26435
rect 15568 26392 15620 26401
rect 17316 26392 17368 26444
rect 18696 26435 18748 26444
rect 18696 26401 18705 26435
rect 18705 26401 18739 26435
rect 18739 26401 18748 26435
rect 18696 26392 18748 26401
rect 19064 26392 19116 26444
rect 21088 26435 21140 26444
rect 21088 26401 21097 26435
rect 21097 26401 21131 26435
rect 21131 26401 21140 26435
rect 21088 26392 21140 26401
rect 22284 26392 22336 26444
rect 26332 26469 26341 26503
rect 26341 26469 26375 26503
rect 26375 26469 26384 26503
rect 26332 26460 26384 26469
rect 30104 26460 30156 26512
rect 25320 26435 25372 26444
rect 7840 26231 7892 26240
rect 7840 26197 7849 26231
rect 7849 26197 7883 26231
rect 7883 26197 7892 26231
rect 7840 26188 7892 26197
rect 9036 26188 9088 26240
rect 11244 26367 11296 26376
rect 11244 26333 11253 26367
rect 11253 26333 11287 26367
rect 11287 26333 11296 26367
rect 11244 26324 11296 26333
rect 11428 26324 11480 26376
rect 20904 26324 20956 26376
rect 22376 26324 22428 26376
rect 11888 26188 11940 26240
rect 12808 26256 12860 26308
rect 18788 26256 18840 26308
rect 25320 26401 25329 26435
rect 25329 26401 25363 26435
rect 25363 26401 25372 26435
rect 25320 26392 25372 26401
rect 25412 26392 25464 26444
rect 33508 26460 33560 26512
rect 31300 26435 31352 26444
rect 24860 26324 24912 26376
rect 27620 26324 27672 26376
rect 31300 26401 31309 26435
rect 31309 26401 31343 26435
rect 31343 26401 31352 26435
rect 31300 26392 31352 26401
rect 30564 26324 30616 26376
rect 32588 26392 32640 26444
rect 33048 26392 33100 26444
rect 31760 26367 31812 26376
rect 31760 26333 31769 26367
rect 31769 26333 31803 26367
rect 31803 26333 31812 26367
rect 31760 26324 31812 26333
rect 24952 26256 25004 26308
rect 25504 26299 25556 26308
rect 25504 26265 25513 26299
rect 25513 26265 25547 26299
rect 25547 26265 25556 26299
rect 25504 26256 25556 26265
rect 12624 26231 12676 26240
rect 12624 26197 12633 26231
rect 12633 26197 12667 26231
rect 12667 26197 12676 26231
rect 12624 26188 12676 26197
rect 29368 26188 29420 26240
rect 31760 26188 31812 26240
rect 6517 26086 6569 26138
rect 6581 26086 6633 26138
rect 6645 26086 6697 26138
rect 6709 26086 6761 26138
rect 17588 26086 17640 26138
rect 17652 26086 17704 26138
rect 17716 26086 17768 26138
rect 17780 26086 17832 26138
rect 28658 26086 28710 26138
rect 28722 26086 28774 26138
rect 28786 26086 28838 26138
rect 28850 26086 28902 26138
rect 5540 25984 5592 26036
rect 8668 25984 8720 26036
rect 10416 25984 10468 26036
rect 13820 25984 13872 26036
rect 14556 26027 14608 26036
rect 14556 25993 14565 26027
rect 14565 25993 14599 26027
rect 14599 25993 14608 26027
rect 14556 25984 14608 25993
rect 15016 25984 15068 26036
rect 7196 25916 7248 25968
rect 9772 25916 9824 25968
rect 3240 25848 3292 25900
rect 7288 25891 7340 25900
rect 5080 25823 5132 25832
rect 5080 25789 5089 25823
rect 5089 25789 5123 25823
rect 5123 25789 5132 25823
rect 5080 25780 5132 25789
rect 5264 25780 5316 25832
rect 2780 25712 2832 25764
rect 4988 25644 5040 25696
rect 7288 25857 7297 25891
rect 7297 25857 7331 25891
rect 7331 25857 7340 25891
rect 7288 25848 7340 25857
rect 7472 25891 7524 25900
rect 7472 25857 7481 25891
rect 7481 25857 7515 25891
rect 7515 25857 7524 25891
rect 7472 25848 7524 25857
rect 9036 25848 9088 25900
rect 7840 25780 7892 25832
rect 7380 25712 7432 25764
rect 8760 25780 8812 25832
rect 10324 25823 10376 25832
rect 10324 25789 10333 25823
rect 10333 25789 10367 25823
rect 10367 25789 10376 25823
rect 10324 25780 10376 25789
rect 11152 25916 11204 25968
rect 11428 25916 11480 25968
rect 12440 25916 12492 25968
rect 20720 25984 20772 26036
rect 22468 25984 22520 26036
rect 26516 25984 26568 26036
rect 27528 25984 27580 26036
rect 30380 25984 30432 26036
rect 30932 25959 30984 25968
rect 13636 25848 13688 25900
rect 20444 25848 20496 25900
rect 26332 25891 26384 25900
rect 11704 25780 11756 25832
rect 10784 25712 10836 25764
rect 11796 25712 11848 25764
rect 12348 25780 12400 25832
rect 15200 25823 15252 25832
rect 15200 25789 15209 25823
rect 15209 25789 15243 25823
rect 15243 25789 15252 25823
rect 15200 25780 15252 25789
rect 16672 25780 16724 25832
rect 17408 25780 17460 25832
rect 17500 25823 17552 25832
rect 17500 25789 17509 25823
rect 17509 25789 17543 25823
rect 17543 25789 17552 25823
rect 17500 25780 17552 25789
rect 19156 25780 19208 25832
rect 23020 25823 23072 25832
rect 23020 25789 23029 25823
rect 23029 25789 23063 25823
rect 23063 25789 23072 25823
rect 23020 25780 23072 25789
rect 13176 25712 13228 25764
rect 14556 25712 14608 25764
rect 15476 25712 15528 25764
rect 20168 25712 20220 25764
rect 23480 25780 23532 25832
rect 26332 25857 26341 25891
rect 26341 25857 26375 25891
rect 26375 25857 26384 25891
rect 26332 25848 26384 25857
rect 26516 25891 26568 25900
rect 26516 25857 26525 25891
rect 26525 25857 26559 25891
rect 26559 25857 26568 25891
rect 26516 25848 26568 25857
rect 23848 25712 23900 25764
rect 24124 25712 24176 25764
rect 25320 25823 25372 25832
rect 25320 25789 25329 25823
rect 25329 25789 25363 25823
rect 25363 25789 25372 25823
rect 25320 25780 25372 25789
rect 24952 25712 25004 25764
rect 25964 25712 26016 25764
rect 7472 25644 7524 25696
rect 9036 25687 9088 25696
rect 9036 25653 9045 25687
rect 9045 25653 9079 25687
rect 9079 25653 9088 25687
rect 9036 25644 9088 25653
rect 9496 25687 9548 25696
rect 9496 25653 9505 25687
rect 9505 25653 9539 25687
rect 9539 25653 9548 25687
rect 9496 25644 9548 25653
rect 11888 25644 11940 25696
rect 12900 25644 12952 25696
rect 16028 25687 16080 25696
rect 16028 25653 16037 25687
rect 16037 25653 16071 25687
rect 16071 25653 16080 25687
rect 16028 25644 16080 25653
rect 16580 25644 16632 25696
rect 23940 25644 23992 25696
rect 25872 25687 25924 25696
rect 25872 25653 25881 25687
rect 25881 25653 25915 25687
rect 25915 25653 25924 25687
rect 25872 25644 25924 25653
rect 30932 25925 30941 25959
rect 30941 25925 30975 25959
rect 30975 25925 30984 25959
rect 30932 25916 30984 25925
rect 28448 25848 28500 25900
rect 26976 25780 27028 25832
rect 30748 25823 30800 25832
rect 30748 25789 30757 25823
rect 30757 25789 30791 25823
rect 30791 25789 30800 25823
rect 30748 25780 30800 25789
rect 31300 25780 31352 25832
rect 31392 25823 31444 25832
rect 31392 25789 31401 25823
rect 31401 25789 31435 25823
rect 31435 25789 31444 25823
rect 33048 25823 33100 25832
rect 31392 25780 31444 25789
rect 33048 25789 33057 25823
rect 33057 25789 33091 25823
rect 33091 25789 33100 25823
rect 33048 25780 33100 25789
rect 33508 25780 33560 25832
rect 28540 25712 28592 25764
rect 29828 25712 29880 25764
rect 31668 25644 31720 25696
rect 12052 25542 12104 25594
rect 12116 25542 12168 25594
rect 12180 25542 12232 25594
rect 12244 25542 12296 25594
rect 23123 25542 23175 25594
rect 23187 25542 23239 25594
rect 23251 25542 23303 25594
rect 23315 25542 23367 25594
rect 1768 25347 1820 25356
rect 1768 25313 1777 25347
rect 1777 25313 1811 25347
rect 1811 25313 1820 25347
rect 1768 25304 1820 25313
rect 2964 25372 3016 25424
rect 3332 25304 3384 25356
rect 5264 25440 5316 25492
rect 8300 25440 8352 25492
rect 12624 25440 12676 25492
rect 13176 25440 13228 25492
rect 5540 25372 5592 25424
rect 7012 25372 7064 25424
rect 9496 25372 9548 25424
rect 12808 25415 12860 25424
rect 12808 25381 12817 25415
rect 12817 25381 12851 25415
rect 12851 25381 12860 25415
rect 12808 25372 12860 25381
rect 18788 25372 18840 25424
rect 23940 25415 23992 25424
rect 2780 25279 2832 25288
rect 2780 25245 2789 25279
rect 2789 25245 2823 25279
rect 2823 25245 2832 25279
rect 2780 25236 2832 25245
rect 2964 25236 3016 25288
rect 4896 25347 4948 25356
rect 4896 25313 4905 25347
rect 4905 25313 4939 25347
rect 4939 25313 4948 25347
rect 4896 25304 4948 25313
rect 7380 25347 7432 25356
rect 7380 25313 7389 25347
rect 7389 25313 7423 25347
rect 7423 25313 7432 25347
rect 7932 25347 7984 25356
rect 7380 25304 7432 25313
rect 7932 25313 7941 25347
rect 7941 25313 7975 25347
rect 7975 25313 7984 25347
rect 7932 25304 7984 25313
rect 9864 25347 9916 25356
rect 9864 25313 9873 25347
rect 9873 25313 9907 25347
rect 9907 25313 9916 25347
rect 9864 25304 9916 25313
rect 10876 25347 10928 25356
rect 10876 25313 10885 25347
rect 10885 25313 10919 25347
rect 10919 25313 10928 25347
rect 10876 25304 10928 25313
rect 11152 25347 11204 25356
rect 11152 25313 11161 25347
rect 11161 25313 11195 25347
rect 11195 25313 11204 25347
rect 11152 25304 11204 25313
rect 11428 25304 11480 25356
rect 12440 25347 12492 25356
rect 12440 25313 12449 25347
rect 12449 25313 12483 25347
rect 12483 25313 12492 25347
rect 12440 25304 12492 25313
rect 12532 25347 12584 25356
rect 12532 25313 12541 25347
rect 12541 25313 12575 25347
rect 12575 25313 12584 25347
rect 12532 25304 12584 25313
rect 5172 25279 5224 25288
rect 5172 25245 5181 25279
rect 5181 25245 5215 25279
rect 5215 25245 5224 25279
rect 5172 25236 5224 25245
rect 7104 25279 7156 25288
rect 7104 25245 7113 25279
rect 7113 25245 7147 25279
rect 7147 25245 7156 25279
rect 7104 25236 7156 25245
rect 7472 25168 7524 25220
rect 2964 25143 3016 25152
rect 2964 25109 2973 25143
rect 2973 25109 3007 25143
rect 3007 25109 3016 25143
rect 2964 25100 3016 25109
rect 4436 25100 4488 25152
rect 5632 25143 5684 25152
rect 5632 25109 5641 25143
rect 5641 25109 5675 25143
rect 5675 25109 5684 25143
rect 5632 25100 5684 25109
rect 9496 25143 9548 25152
rect 9496 25109 9505 25143
rect 9505 25109 9539 25143
rect 9539 25109 9548 25143
rect 9496 25100 9548 25109
rect 10048 25168 10100 25220
rect 12164 25168 12216 25220
rect 12900 25347 12952 25356
rect 12900 25313 12909 25347
rect 12909 25313 12943 25347
rect 12943 25313 12952 25347
rect 12900 25304 12952 25313
rect 16212 25304 16264 25356
rect 18144 25304 18196 25356
rect 22928 25304 22980 25356
rect 23480 25347 23532 25356
rect 23480 25313 23489 25347
rect 23489 25313 23523 25347
rect 23523 25313 23532 25347
rect 23480 25304 23532 25313
rect 23940 25381 23949 25415
rect 23949 25381 23983 25415
rect 23983 25381 23992 25415
rect 23940 25372 23992 25381
rect 24124 25347 24176 25356
rect 24124 25313 24133 25347
rect 24133 25313 24167 25347
rect 24167 25313 24176 25347
rect 24124 25304 24176 25313
rect 13820 25236 13872 25288
rect 14924 25236 14976 25288
rect 19156 25236 19208 25288
rect 13728 25168 13780 25220
rect 17500 25168 17552 25220
rect 16672 25100 16724 25152
rect 17132 25100 17184 25152
rect 23848 25100 23900 25152
rect 25320 25440 25372 25492
rect 28540 25483 28592 25492
rect 28540 25449 28549 25483
rect 28549 25449 28583 25483
rect 28583 25449 28592 25483
rect 28540 25440 28592 25449
rect 31392 25440 31444 25492
rect 25872 25372 25924 25424
rect 28172 25347 28224 25356
rect 28172 25313 28181 25347
rect 28181 25313 28215 25347
rect 28215 25313 28224 25347
rect 28172 25304 28224 25313
rect 28448 25304 28500 25356
rect 29368 25347 29420 25356
rect 29368 25313 29377 25347
rect 29377 25313 29411 25347
rect 29411 25313 29420 25347
rect 29368 25304 29420 25313
rect 31668 25372 31720 25424
rect 31576 25347 31628 25356
rect 26884 25236 26936 25288
rect 31576 25313 31585 25347
rect 31585 25313 31619 25347
rect 31619 25313 31628 25347
rect 31576 25304 31628 25313
rect 31760 25347 31812 25356
rect 31760 25313 31769 25347
rect 31769 25313 31803 25347
rect 31803 25313 31812 25347
rect 31760 25304 31812 25313
rect 33324 25304 33376 25356
rect 33508 25347 33560 25356
rect 33508 25313 33517 25347
rect 33517 25313 33551 25347
rect 33551 25313 33560 25347
rect 33508 25304 33560 25313
rect 31852 25168 31904 25220
rect 33140 25100 33192 25152
rect 6517 24998 6569 25050
rect 6581 24998 6633 25050
rect 6645 24998 6697 25050
rect 6709 24998 6761 25050
rect 17588 24998 17640 25050
rect 17652 24998 17704 25050
rect 17716 24998 17768 25050
rect 17780 24998 17832 25050
rect 28658 24998 28710 25050
rect 28722 24998 28774 25050
rect 28786 24998 28838 25050
rect 28850 24998 28902 25050
rect 4896 24896 4948 24948
rect 7104 24896 7156 24948
rect 7288 24896 7340 24948
rect 5080 24760 5132 24812
rect 1492 24692 1544 24744
rect 2964 24624 3016 24676
rect 4436 24735 4488 24744
rect 5632 24760 5684 24812
rect 9588 24828 9640 24880
rect 9772 24896 9824 24948
rect 10232 24896 10284 24948
rect 15016 24896 15068 24948
rect 16212 24939 16264 24948
rect 16212 24905 16221 24939
rect 16221 24905 16255 24939
rect 16255 24905 16264 24939
rect 16212 24896 16264 24905
rect 30748 24939 30800 24948
rect 30748 24905 30757 24939
rect 30757 24905 30791 24939
rect 30791 24905 30800 24939
rect 30748 24896 30800 24905
rect 12164 24828 12216 24880
rect 14004 24828 14056 24880
rect 14924 24828 14976 24880
rect 10784 24803 10836 24812
rect 10784 24769 10793 24803
rect 10793 24769 10827 24803
rect 10827 24769 10836 24803
rect 10784 24760 10836 24769
rect 11888 24760 11940 24812
rect 16304 24803 16356 24812
rect 4436 24701 4454 24735
rect 4454 24701 4488 24735
rect 4436 24692 4488 24701
rect 7196 24735 7248 24744
rect 7196 24701 7205 24735
rect 7205 24701 7239 24735
rect 7239 24701 7248 24735
rect 7196 24692 7248 24701
rect 8300 24735 8352 24744
rect 8300 24701 8309 24735
rect 8309 24701 8343 24735
rect 8343 24701 8352 24735
rect 8300 24692 8352 24701
rect 9496 24692 9548 24744
rect 10232 24735 10284 24744
rect 10232 24701 10241 24735
rect 10241 24701 10275 24735
rect 10275 24701 10284 24735
rect 10232 24692 10284 24701
rect 12256 24735 12308 24744
rect 5080 24624 5132 24676
rect 9404 24624 9456 24676
rect 9956 24624 10008 24676
rect 12256 24701 12265 24735
rect 12265 24701 12299 24735
rect 12299 24701 12308 24735
rect 12256 24692 12308 24701
rect 12992 24692 13044 24744
rect 13636 24735 13688 24744
rect 13636 24701 13645 24735
rect 13645 24701 13679 24735
rect 13679 24701 13688 24735
rect 13636 24692 13688 24701
rect 15292 24735 15344 24744
rect 15292 24701 15301 24735
rect 15301 24701 15335 24735
rect 15335 24701 15344 24735
rect 15292 24692 15344 24701
rect 16028 24735 16080 24744
rect 16028 24701 16037 24735
rect 16037 24701 16071 24735
rect 16071 24701 16080 24735
rect 16028 24692 16080 24701
rect 16304 24769 16313 24803
rect 16313 24769 16347 24803
rect 16347 24769 16356 24803
rect 16304 24760 16356 24769
rect 16672 24760 16724 24812
rect 16580 24692 16632 24744
rect 17408 24692 17460 24744
rect 19156 24760 19208 24812
rect 20168 24760 20220 24812
rect 13360 24624 13412 24676
rect 14372 24624 14424 24676
rect 15200 24624 15252 24676
rect 17132 24624 17184 24676
rect 19432 24624 19484 24676
rect 2136 24556 2188 24608
rect 3332 24599 3384 24608
rect 3332 24565 3341 24599
rect 3341 24565 3375 24599
rect 3375 24565 3384 24599
rect 3332 24556 3384 24565
rect 5172 24556 5224 24608
rect 8852 24599 8904 24608
rect 8852 24565 8861 24599
rect 8861 24565 8895 24599
rect 8895 24565 8904 24599
rect 8852 24556 8904 24565
rect 9864 24556 9916 24608
rect 11244 24556 11296 24608
rect 13820 24599 13872 24608
rect 13820 24565 13829 24599
rect 13829 24565 13863 24599
rect 13863 24565 13872 24599
rect 13820 24556 13872 24565
rect 17224 24556 17276 24608
rect 19524 24556 19576 24608
rect 21088 24692 21140 24744
rect 22928 24760 22980 24812
rect 23480 24803 23532 24812
rect 23480 24769 23489 24803
rect 23489 24769 23523 24803
rect 23523 24769 23532 24803
rect 23480 24760 23532 24769
rect 20444 24624 20496 24676
rect 23020 24624 23072 24676
rect 20536 24556 20588 24608
rect 20812 24556 20864 24608
rect 22560 24556 22612 24608
rect 23756 24735 23808 24744
rect 23756 24701 23765 24735
rect 23765 24701 23799 24735
rect 23799 24701 23808 24735
rect 23756 24692 23808 24701
rect 23940 24692 23992 24744
rect 25044 24735 25096 24744
rect 25044 24701 25053 24735
rect 25053 24701 25087 24735
rect 25087 24701 25096 24735
rect 25044 24692 25096 24701
rect 28172 24692 28224 24744
rect 29184 24692 29236 24744
rect 30472 24760 30524 24812
rect 30932 24760 30984 24812
rect 33324 24803 33376 24812
rect 33324 24769 33333 24803
rect 33333 24769 33367 24803
rect 33367 24769 33376 24803
rect 33324 24760 33376 24769
rect 23848 24624 23900 24676
rect 26424 24624 26476 24676
rect 30748 24692 30800 24744
rect 32128 24735 32180 24744
rect 32128 24701 32137 24735
rect 32137 24701 32171 24735
rect 32171 24701 32180 24735
rect 32128 24692 32180 24701
rect 32956 24692 33008 24744
rect 33232 24735 33284 24744
rect 33232 24701 33241 24735
rect 33241 24701 33275 24735
rect 33275 24701 33284 24735
rect 33232 24692 33284 24701
rect 31760 24624 31812 24676
rect 25228 24599 25280 24608
rect 25228 24565 25237 24599
rect 25237 24565 25271 24599
rect 25271 24565 25280 24599
rect 25228 24556 25280 24565
rect 27160 24556 27212 24608
rect 28264 24556 28316 24608
rect 28356 24556 28408 24608
rect 12052 24454 12104 24506
rect 12116 24454 12168 24506
rect 12180 24454 12232 24506
rect 12244 24454 12296 24506
rect 23123 24454 23175 24506
rect 23187 24454 23239 24506
rect 23251 24454 23303 24506
rect 23315 24454 23367 24506
rect 7564 24352 7616 24404
rect 2872 24284 2924 24336
rect 6276 24327 6328 24336
rect 6276 24293 6285 24327
rect 6285 24293 6319 24327
rect 6319 24293 6328 24327
rect 9036 24352 9088 24404
rect 10600 24352 10652 24404
rect 6276 24284 6328 24293
rect 7932 24284 7984 24336
rect 10784 24284 10836 24336
rect 11244 24327 11296 24336
rect 11244 24293 11253 24327
rect 11253 24293 11287 24327
rect 11287 24293 11296 24327
rect 11244 24284 11296 24293
rect 11612 24352 11664 24404
rect 1400 24259 1452 24268
rect 1400 24225 1409 24259
rect 1409 24225 1443 24259
rect 1443 24225 1452 24259
rect 1400 24216 1452 24225
rect 2136 24259 2188 24268
rect 2136 24225 2145 24259
rect 2145 24225 2179 24259
rect 2179 24225 2188 24259
rect 2136 24216 2188 24225
rect 3332 24259 3384 24268
rect 3332 24225 3341 24259
rect 3341 24225 3375 24259
rect 3375 24225 3384 24259
rect 3332 24216 3384 24225
rect 4344 24216 4396 24268
rect 5172 24259 5224 24268
rect 5172 24225 5181 24259
rect 5181 24225 5215 24259
rect 5215 24225 5224 24259
rect 5172 24216 5224 24225
rect 6920 24216 6972 24268
rect 4528 24148 4580 24200
rect 3792 24080 3844 24132
rect 4620 24123 4672 24132
rect 4620 24089 4629 24123
rect 4629 24089 4663 24123
rect 4663 24089 4672 24123
rect 4620 24080 4672 24089
rect 1768 24012 1820 24064
rect 2780 24012 2832 24064
rect 7564 24216 7616 24268
rect 11796 24216 11848 24268
rect 11244 24148 11296 24200
rect 11520 24191 11572 24200
rect 11520 24157 11529 24191
rect 11529 24157 11563 24191
rect 11563 24157 11572 24191
rect 11520 24148 11572 24157
rect 12348 24148 12400 24200
rect 12992 24395 13044 24404
rect 12992 24361 13001 24395
rect 13001 24361 13035 24395
rect 13035 24361 13044 24395
rect 18144 24395 18196 24404
rect 12992 24352 13044 24361
rect 18144 24361 18153 24395
rect 18153 24361 18187 24395
rect 18187 24361 18196 24395
rect 18144 24352 18196 24361
rect 16304 24284 16356 24336
rect 17132 24259 17184 24268
rect 14556 24148 14608 24200
rect 17132 24225 17141 24259
rect 17141 24225 17175 24259
rect 17175 24225 17184 24259
rect 17132 24216 17184 24225
rect 17224 24191 17276 24200
rect 17224 24157 17233 24191
rect 17233 24157 17267 24191
rect 17267 24157 17276 24191
rect 17224 24148 17276 24157
rect 8668 24080 8720 24132
rect 9956 24080 10008 24132
rect 11704 24080 11756 24132
rect 15292 24080 15344 24132
rect 16120 24123 16172 24132
rect 16120 24089 16129 24123
rect 16129 24089 16163 24123
rect 16163 24089 16172 24123
rect 16120 24080 16172 24089
rect 20444 24352 20496 24404
rect 21088 24352 21140 24404
rect 22928 24352 22980 24404
rect 25136 24352 25188 24404
rect 18788 24284 18840 24336
rect 22376 24284 22428 24336
rect 23020 24284 23072 24336
rect 20996 24191 21048 24200
rect 20996 24157 21005 24191
rect 21005 24157 21039 24191
rect 21039 24157 21048 24191
rect 20996 24148 21048 24157
rect 21364 24191 21416 24200
rect 21364 24157 21373 24191
rect 21373 24157 21407 24191
rect 21407 24157 21416 24191
rect 21364 24148 21416 24157
rect 23940 24284 23992 24336
rect 23848 24216 23900 24268
rect 27896 24352 27948 24404
rect 29184 24395 29236 24404
rect 29184 24361 29193 24395
rect 29193 24361 29227 24395
rect 29227 24361 29236 24395
rect 29184 24352 29236 24361
rect 31208 24395 31260 24404
rect 31208 24361 31217 24395
rect 31217 24361 31251 24395
rect 31251 24361 31260 24395
rect 31208 24352 31260 24361
rect 27160 24327 27212 24336
rect 27160 24293 27169 24327
rect 27169 24293 27203 24327
rect 27203 24293 27212 24327
rect 27160 24284 27212 24293
rect 28448 24284 28500 24336
rect 25504 24259 25556 24268
rect 25504 24225 25513 24259
rect 25513 24225 25547 24259
rect 25547 24225 25556 24259
rect 25504 24216 25556 24225
rect 25872 24259 25924 24268
rect 25872 24225 25881 24259
rect 25881 24225 25915 24259
rect 25915 24225 25924 24259
rect 25872 24216 25924 24225
rect 25964 24259 26016 24268
rect 25964 24225 25973 24259
rect 25973 24225 26007 24259
rect 26007 24225 26016 24259
rect 25964 24216 26016 24225
rect 26884 24191 26936 24200
rect 26884 24157 26893 24191
rect 26893 24157 26927 24191
rect 26927 24157 26936 24191
rect 26884 24148 26936 24157
rect 28356 24148 28408 24200
rect 28540 24148 28592 24200
rect 30840 24216 30892 24268
rect 31392 24148 31444 24200
rect 31760 24148 31812 24200
rect 32128 24284 32180 24336
rect 32588 24284 32640 24336
rect 32864 24148 32916 24200
rect 11612 24012 11664 24064
rect 12256 24055 12308 24064
rect 12256 24021 12265 24055
rect 12265 24021 12299 24055
rect 12299 24021 12308 24055
rect 12256 24012 12308 24021
rect 12900 24012 12952 24064
rect 17960 24012 18012 24064
rect 23020 24012 23072 24064
rect 29828 24080 29880 24132
rect 23664 24055 23716 24064
rect 23664 24021 23673 24055
rect 23673 24021 23707 24055
rect 23707 24021 23716 24055
rect 23664 24012 23716 24021
rect 24400 24012 24452 24064
rect 30748 24055 30800 24064
rect 30748 24021 30757 24055
rect 30757 24021 30791 24055
rect 30791 24021 30800 24055
rect 30748 24012 30800 24021
rect 33600 24055 33652 24064
rect 33600 24021 33609 24055
rect 33609 24021 33643 24055
rect 33643 24021 33652 24055
rect 33600 24012 33652 24021
rect 6517 23910 6569 23962
rect 6581 23910 6633 23962
rect 6645 23910 6697 23962
rect 6709 23910 6761 23962
rect 17588 23910 17640 23962
rect 17652 23910 17704 23962
rect 17716 23910 17768 23962
rect 17780 23910 17832 23962
rect 28658 23910 28710 23962
rect 28722 23910 28774 23962
rect 28786 23910 28838 23962
rect 28850 23910 28902 23962
rect 2964 23808 3016 23860
rect 8852 23808 8904 23860
rect 9588 23808 9640 23860
rect 10600 23808 10652 23860
rect 11704 23808 11756 23860
rect 12348 23851 12400 23860
rect 12348 23817 12357 23851
rect 12357 23817 12391 23851
rect 12391 23817 12400 23851
rect 12348 23808 12400 23817
rect 19432 23851 19484 23860
rect 19432 23817 19441 23851
rect 19441 23817 19475 23851
rect 19475 23817 19484 23851
rect 19432 23808 19484 23817
rect 26884 23808 26936 23860
rect 4344 23740 4396 23792
rect 4436 23715 4488 23724
rect 4436 23681 4445 23715
rect 4445 23681 4479 23715
rect 4479 23681 4488 23715
rect 4436 23672 4488 23681
rect 4620 23672 4672 23724
rect 11520 23740 11572 23792
rect 29460 23783 29512 23792
rect 4896 23604 4948 23656
rect 5264 23604 5316 23656
rect 6920 23604 6972 23656
rect 9128 23672 9180 23724
rect 3332 23579 3384 23588
rect 3332 23545 3341 23579
rect 3341 23545 3375 23579
rect 3375 23545 3384 23579
rect 3332 23536 3384 23545
rect 9220 23604 9272 23656
rect 10232 23672 10284 23724
rect 10324 23672 10376 23724
rect 9772 23647 9824 23656
rect 9772 23613 9781 23647
rect 9781 23613 9815 23647
rect 9815 23613 9824 23647
rect 9772 23604 9824 23613
rect 9956 23647 10008 23656
rect 9956 23613 9965 23647
rect 9965 23613 9999 23647
rect 9999 23613 10008 23647
rect 9956 23604 10008 23613
rect 8392 23468 8444 23520
rect 8484 23468 8536 23520
rect 11428 23604 11480 23656
rect 12440 23672 12492 23724
rect 29460 23749 29469 23783
rect 29469 23749 29503 23783
rect 29503 23749 29512 23783
rect 29460 23740 29512 23749
rect 12900 23672 12952 23724
rect 12624 23536 12676 23588
rect 14556 23604 14608 23656
rect 15476 23604 15528 23656
rect 13728 23536 13780 23588
rect 20628 23536 20680 23588
rect 23480 23604 23532 23656
rect 23848 23647 23900 23656
rect 23848 23613 23857 23647
rect 23857 23613 23891 23647
rect 23891 23613 23900 23647
rect 23848 23604 23900 23613
rect 24400 23604 24452 23656
rect 25228 23672 25280 23724
rect 28448 23672 28500 23724
rect 30748 23672 30800 23724
rect 28540 23647 28592 23656
rect 23572 23536 23624 23588
rect 24308 23579 24360 23588
rect 24308 23545 24317 23579
rect 24317 23545 24351 23579
rect 24351 23545 24360 23579
rect 24308 23536 24360 23545
rect 24492 23536 24544 23588
rect 28540 23613 28549 23647
rect 28549 23613 28583 23647
rect 28583 23613 28592 23647
rect 28540 23604 28592 23613
rect 29644 23647 29696 23656
rect 29644 23613 29653 23647
rect 29653 23613 29687 23647
rect 29687 23613 29696 23647
rect 29644 23604 29696 23613
rect 30472 23647 30524 23656
rect 30472 23613 30481 23647
rect 30481 23613 30515 23647
rect 30515 23613 30524 23647
rect 30472 23604 30524 23613
rect 31852 23647 31904 23656
rect 31852 23613 31861 23647
rect 31861 23613 31895 23647
rect 31895 23613 31904 23647
rect 31852 23604 31904 23613
rect 25504 23536 25556 23588
rect 13268 23468 13320 23520
rect 13636 23468 13688 23520
rect 19616 23511 19668 23520
rect 19616 23477 19625 23511
rect 19625 23477 19659 23511
rect 19659 23477 19668 23511
rect 19616 23468 19668 23477
rect 20168 23468 20220 23520
rect 20996 23468 21048 23520
rect 26792 23511 26844 23520
rect 26792 23477 26801 23511
rect 26801 23477 26835 23511
rect 26835 23477 26844 23511
rect 26792 23468 26844 23477
rect 28172 23511 28224 23520
rect 28172 23477 28181 23511
rect 28181 23477 28215 23511
rect 28215 23477 28224 23511
rect 28172 23468 28224 23477
rect 30656 23536 30708 23588
rect 12052 23366 12104 23418
rect 12116 23366 12168 23418
rect 12180 23366 12232 23418
rect 12244 23366 12296 23418
rect 23123 23366 23175 23418
rect 23187 23366 23239 23418
rect 23251 23366 23303 23418
rect 23315 23366 23367 23418
rect 9128 23264 9180 23316
rect 9956 23264 10008 23316
rect 2688 23196 2740 23248
rect 5172 23196 5224 23248
rect 2964 23128 3016 23180
rect 7104 23171 7156 23180
rect 7104 23137 7113 23171
rect 7113 23137 7147 23171
rect 7147 23137 7156 23171
rect 7104 23128 7156 23137
rect 9772 23196 9824 23248
rect 10048 23171 10100 23180
rect 10048 23137 10057 23171
rect 10057 23137 10091 23171
rect 10091 23137 10100 23171
rect 10048 23128 10100 23137
rect 11060 23264 11112 23316
rect 11888 23264 11940 23316
rect 14188 23264 14240 23316
rect 14740 23264 14792 23316
rect 17408 23264 17460 23316
rect 11428 23196 11480 23248
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 4160 23060 4212 23112
rect 5356 23103 5408 23112
rect 5356 23069 5365 23103
rect 5365 23069 5399 23103
rect 5399 23069 5408 23103
rect 5356 23060 5408 23069
rect 5816 23060 5868 23112
rect 9312 23060 9364 23112
rect 11244 23128 11296 23180
rect 12440 23196 12492 23248
rect 16120 23239 16172 23248
rect 16120 23205 16154 23239
rect 16154 23205 16172 23239
rect 16120 23196 16172 23205
rect 16304 23196 16356 23248
rect 16672 23196 16724 23248
rect 17960 23264 18012 23316
rect 21364 23264 21416 23316
rect 25504 23264 25556 23316
rect 19616 23196 19668 23248
rect 23020 23196 23072 23248
rect 23480 23196 23532 23248
rect 24400 23196 24452 23248
rect 25136 23196 25188 23248
rect 28448 23264 28500 23316
rect 26792 23196 26844 23248
rect 28264 23196 28316 23248
rect 12716 23128 12768 23180
rect 15016 23128 15068 23180
rect 17224 23128 17276 23180
rect 18696 23128 18748 23180
rect 14372 23060 14424 23112
rect 19340 23128 19392 23180
rect 19524 23060 19576 23112
rect 20444 23128 20496 23180
rect 20720 23171 20772 23180
rect 20720 23137 20729 23171
rect 20729 23137 20763 23171
rect 20763 23137 20772 23171
rect 22376 23171 22428 23180
rect 20720 23128 20772 23137
rect 22376 23137 22385 23171
rect 22385 23137 22419 23171
rect 22419 23137 22428 23171
rect 22376 23128 22428 23137
rect 24768 23128 24820 23180
rect 25964 23128 26016 23180
rect 28172 23128 28224 23180
rect 20812 23060 20864 23112
rect 21732 23103 21784 23112
rect 21732 23069 21741 23103
rect 21741 23069 21775 23103
rect 21775 23069 21784 23103
rect 21732 23060 21784 23069
rect 25780 23060 25832 23112
rect 29368 23128 29420 23180
rect 31760 23264 31812 23316
rect 32864 23307 32916 23316
rect 32864 23273 32873 23307
rect 32873 23273 32907 23307
rect 32907 23273 32916 23307
rect 32864 23264 32916 23273
rect 32956 23264 33008 23316
rect 33600 23264 33652 23316
rect 32588 23128 32640 23180
rect 30932 23103 30984 23112
rect 4896 22992 4948 23044
rect 8024 23035 8076 23044
rect 8024 23001 8033 23035
rect 8033 23001 8067 23035
rect 8067 23001 8076 23035
rect 8024 22992 8076 23001
rect 8300 22992 8352 23044
rect 10876 22992 10928 23044
rect 4712 22924 4764 22976
rect 12992 22924 13044 22976
rect 18788 22967 18840 22976
rect 18788 22933 18797 22967
rect 18797 22933 18831 22967
rect 18831 22933 18840 22967
rect 18788 22924 18840 22933
rect 23480 22924 23532 22976
rect 23848 22992 23900 23044
rect 27804 22992 27856 23044
rect 30932 23069 30941 23103
rect 30941 23069 30975 23103
rect 30975 23069 30984 23103
rect 30932 23060 30984 23069
rect 31024 23060 31076 23112
rect 30012 22992 30064 23044
rect 27528 22924 27580 22976
rect 28540 22924 28592 22976
rect 31392 22924 31444 22976
rect 6517 22822 6569 22874
rect 6581 22822 6633 22874
rect 6645 22822 6697 22874
rect 6709 22822 6761 22874
rect 17588 22822 17640 22874
rect 17652 22822 17704 22874
rect 17716 22822 17768 22874
rect 17780 22822 17832 22874
rect 28658 22822 28710 22874
rect 28722 22822 28774 22874
rect 28786 22822 28838 22874
rect 28850 22822 28902 22874
rect 3332 22720 3384 22772
rect 4160 22763 4212 22772
rect 4160 22729 4169 22763
rect 4169 22729 4203 22763
rect 4203 22729 4212 22763
rect 4160 22720 4212 22729
rect 6920 22763 6972 22772
rect 6920 22729 6929 22763
rect 6929 22729 6963 22763
rect 6963 22729 6972 22763
rect 6920 22720 6972 22729
rect 10232 22720 10284 22772
rect 10968 22763 11020 22772
rect 10968 22729 10977 22763
rect 10977 22729 11011 22763
rect 11011 22729 11020 22763
rect 10968 22720 11020 22729
rect 12992 22763 13044 22772
rect 2688 22652 2740 22704
rect 5816 22695 5868 22704
rect 4712 22584 4764 22636
rect 5816 22661 5825 22695
rect 5825 22661 5859 22695
rect 5859 22661 5868 22695
rect 5816 22652 5868 22661
rect 2688 22559 2740 22568
rect 2688 22525 2697 22559
rect 2697 22525 2731 22559
rect 2731 22525 2740 22559
rect 2688 22516 2740 22525
rect 2964 22516 3016 22568
rect 3332 22559 3384 22568
rect 3332 22525 3341 22559
rect 3341 22525 3375 22559
rect 3375 22525 3384 22559
rect 3332 22516 3384 22525
rect 4344 22559 4396 22568
rect 2780 22423 2832 22432
rect 2780 22389 2789 22423
rect 2789 22389 2823 22423
rect 2823 22389 2832 22423
rect 4344 22525 4353 22559
rect 4353 22525 4387 22559
rect 4387 22525 4396 22559
rect 4344 22516 4396 22525
rect 4436 22559 4488 22568
rect 4436 22525 4445 22559
rect 4445 22525 4479 22559
rect 4479 22525 4488 22559
rect 7012 22584 7064 22636
rect 4436 22516 4488 22525
rect 6276 22516 6328 22568
rect 7932 22584 7984 22636
rect 8392 22627 8444 22636
rect 8392 22593 8401 22627
rect 8401 22593 8435 22627
rect 8435 22593 8444 22627
rect 8392 22584 8444 22593
rect 8760 22584 8812 22636
rect 4712 22491 4764 22500
rect 4712 22457 4721 22491
rect 4721 22457 4755 22491
rect 4755 22457 4764 22491
rect 4712 22448 4764 22457
rect 11152 22516 11204 22568
rect 12992 22729 13001 22763
rect 13001 22729 13035 22763
rect 13035 22729 13044 22763
rect 12992 22720 13044 22729
rect 15016 22720 15068 22772
rect 15568 22720 15620 22772
rect 19524 22763 19576 22772
rect 19524 22729 19533 22763
rect 19533 22729 19567 22763
rect 19567 22729 19576 22763
rect 19524 22720 19576 22729
rect 28264 22720 28316 22772
rect 12532 22652 12584 22704
rect 19616 22652 19668 22704
rect 21824 22652 21876 22704
rect 13176 22627 13228 22636
rect 13176 22593 13185 22627
rect 13185 22593 13219 22627
rect 13219 22593 13228 22627
rect 13176 22584 13228 22593
rect 13820 22584 13872 22636
rect 16304 22584 16356 22636
rect 18788 22627 18840 22636
rect 18788 22593 18797 22627
rect 18797 22593 18831 22627
rect 18831 22593 18840 22627
rect 18788 22584 18840 22593
rect 10968 22448 11020 22500
rect 13360 22516 13412 22568
rect 15476 22516 15528 22568
rect 19432 22516 19484 22568
rect 14372 22491 14424 22500
rect 14372 22457 14381 22491
rect 14381 22457 14415 22491
rect 14415 22457 14424 22491
rect 14372 22448 14424 22457
rect 19340 22448 19392 22500
rect 2780 22380 2832 22389
rect 6736 22380 6788 22432
rect 8024 22380 8076 22432
rect 9312 22423 9364 22432
rect 9312 22389 9321 22423
rect 9321 22389 9355 22423
rect 9355 22389 9364 22423
rect 9312 22380 9364 22389
rect 11796 22380 11848 22432
rect 17316 22423 17368 22432
rect 17316 22389 17325 22423
rect 17325 22389 17359 22423
rect 17359 22389 17368 22423
rect 19984 22516 20036 22568
rect 19708 22448 19760 22500
rect 20536 22448 20588 22500
rect 23572 22652 23624 22704
rect 29828 22720 29880 22772
rect 30012 22763 30064 22772
rect 30012 22729 30021 22763
rect 30021 22729 30055 22763
rect 30055 22729 30064 22763
rect 30012 22720 30064 22729
rect 30932 22720 30984 22772
rect 24768 22584 24820 22636
rect 17316 22380 17368 22389
rect 19892 22380 19944 22432
rect 20352 22380 20404 22432
rect 20628 22423 20680 22432
rect 20628 22389 20637 22423
rect 20637 22389 20671 22423
rect 20671 22389 20680 22423
rect 20628 22380 20680 22389
rect 23020 22516 23072 22568
rect 23664 22516 23716 22568
rect 23848 22559 23900 22568
rect 23848 22525 23857 22559
rect 23857 22525 23891 22559
rect 23891 22525 23900 22559
rect 23848 22516 23900 22525
rect 24032 22516 24084 22568
rect 24400 22559 24452 22568
rect 24400 22525 24409 22559
rect 24409 22525 24443 22559
rect 24443 22525 24452 22559
rect 24400 22516 24452 22525
rect 27068 22584 27120 22636
rect 27528 22584 27580 22636
rect 28540 22627 28592 22636
rect 28540 22593 28549 22627
rect 28549 22593 28583 22627
rect 28583 22593 28592 22627
rect 28540 22584 28592 22593
rect 30840 22584 30892 22636
rect 31392 22627 31444 22636
rect 26884 22516 26936 22568
rect 31392 22593 31401 22627
rect 31401 22593 31435 22627
rect 31435 22593 31444 22627
rect 31392 22584 31444 22593
rect 23940 22380 23992 22432
rect 26148 22423 26200 22432
rect 26148 22389 26157 22423
rect 26157 22389 26191 22423
rect 26191 22389 26200 22423
rect 26148 22380 26200 22389
rect 29828 22448 29880 22500
rect 32588 22448 32640 22500
rect 29368 22380 29420 22432
rect 30932 22380 30984 22432
rect 12052 22278 12104 22330
rect 12116 22278 12168 22330
rect 12180 22278 12232 22330
rect 12244 22278 12296 22330
rect 23123 22278 23175 22330
rect 23187 22278 23239 22330
rect 23251 22278 23303 22330
rect 23315 22278 23367 22330
rect 4712 22176 4764 22228
rect 10324 22176 10376 22228
rect 10876 22176 10928 22228
rect 11704 22176 11756 22228
rect 12348 22219 12400 22228
rect 12348 22185 12357 22219
rect 12357 22185 12391 22219
rect 12391 22185 12400 22219
rect 12348 22176 12400 22185
rect 16580 22176 16632 22228
rect 21456 22176 21508 22228
rect 2688 22108 2740 22160
rect 3332 22108 3384 22160
rect 4252 22108 4304 22160
rect 4620 22040 4672 22092
rect 4896 22083 4948 22092
rect 4896 22049 4905 22083
rect 4905 22049 4939 22083
rect 4939 22049 4948 22083
rect 4896 22040 4948 22049
rect 5356 22083 5408 22092
rect 5356 22049 5365 22083
rect 5365 22049 5399 22083
rect 5399 22049 5408 22083
rect 5356 22040 5408 22049
rect 5540 22083 5592 22092
rect 5540 22049 5549 22083
rect 5549 22049 5583 22083
rect 5583 22049 5592 22083
rect 5540 22040 5592 22049
rect 6736 22108 6788 22160
rect 6920 22083 6972 22092
rect 6920 22049 6929 22083
rect 6929 22049 6963 22083
rect 6963 22049 6972 22083
rect 6920 22040 6972 22049
rect 9312 22108 9364 22160
rect 11060 22108 11112 22160
rect 13820 22108 13872 22160
rect 7472 22040 7524 22092
rect 7932 22040 7984 22092
rect 10784 22040 10836 22092
rect 11152 22083 11204 22092
rect 11152 22049 11161 22083
rect 11161 22049 11195 22083
rect 11195 22049 11204 22083
rect 11152 22040 11204 22049
rect 12348 22083 12400 22092
rect 12348 22049 12357 22083
rect 12357 22049 12391 22083
rect 12391 22049 12400 22083
rect 12348 22040 12400 22049
rect 13360 22083 13412 22092
rect 13360 22049 13369 22083
rect 13369 22049 13403 22083
rect 13403 22049 13412 22083
rect 13360 22040 13412 22049
rect 2780 21972 2832 22024
rect 4068 21972 4120 22024
rect 7104 22015 7156 22024
rect 7104 21981 7113 22015
rect 7113 21981 7147 22015
rect 7147 21981 7156 22015
rect 7104 21972 7156 21981
rect 11888 21972 11940 22024
rect 12532 22015 12584 22024
rect 12532 21981 12541 22015
rect 12541 21981 12575 22015
rect 12575 21981 12584 22015
rect 12532 21972 12584 21981
rect 15292 22040 15344 22092
rect 18604 22108 18656 22160
rect 21732 22108 21784 22160
rect 21824 22108 21876 22160
rect 16580 22083 16632 22092
rect 16580 22049 16589 22083
rect 16589 22049 16623 22083
rect 16623 22049 16632 22083
rect 16580 22040 16632 22049
rect 22744 22083 22796 22092
rect 22744 22049 22753 22083
rect 22753 22049 22787 22083
rect 22787 22049 22796 22083
rect 22744 22040 22796 22049
rect 23572 22040 23624 22092
rect 24400 22040 24452 22092
rect 25780 22040 25832 22092
rect 26148 22040 26200 22092
rect 27068 22083 27120 22092
rect 19432 21972 19484 22024
rect 20168 22015 20220 22024
rect 20168 21981 20177 22015
rect 20177 21981 20211 22015
rect 20211 21981 20220 22015
rect 20168 21972 20220 21981
rect 22376 21972 22428 22024
rect 7288 21904 7340 21956
rect 12164 21904 12216 21956
rect 1676 21836 1728 21888
rect 2964 21836 3016 21888
rect 4988 21836 5040 21888
rect 11244 21836 11296 21888
rect 21824 21904 21876 21956
rect 23940 21972 23992 22024
rect 24492 21972 24544 22024
rect 24768 21972 24820 22024
rect 27068 22049 27077 22083
rect 27077 22049 27111 22083
rect 27111 22049 27120 22083
rect 27068 22040 27120 22049
rect 27436 22083 27488 22092
rect 27436 22049 27445 22083
rect 27445 22049 27479 22083
rect 27479 22049 27488 22083
rect 27436 22040 27488 22049
rect 28172 22108 28224 22160
rect 30840 22151 30892 22160
rect 30840 22117 30870 22151
rect 30870 22117 30892 22151
rect 30840 22108 30892 22117
rect 31852 22108 31904 22160
rect 32036 22083 32088 22092
rect 27988 21972 28040 22024
rect 30656 21904 30708 21956
rect 32036 22049 32045 22083
rect 32045 22049 32079 22083
rect 32079 22049 32088 22083
rect 32036 22040 32088 22049
rect 33048 22040 33100 22092
rect 14832 21836 14884 21888
rect 21916 21879 21968 21888
rect 21916 21845 21925 21879
rect 21925 21845 21959 21879
rect 21959 21845 21968 21879
rect 21916 21836 21968 21845
rect 26516 21836 26568 21888
rect 29644 21836 29696 21888
rect 30932 21836 30984 21888
rect 6517 21734 6569 21786
rect 6581 21734 6633 21786
rect 6645 21734 6697 21786
rect 6709 21734 6761 21786
rect 17588 21734 17640 21786
rect 17652 21734 17704 21786
rect 17716 21734 17768 21786
rect 17780 21734 17832 21786
rect 28658 21734 28710 21786
rect 28722 21734 28774 21786
rect 28786 21734 28838 21786
rect 28850 21734 28902 21786
rect 11152 21675 11204 21684
rect 11152 21641 11161 21675
rect 11161 21641 11195 21675
rect 11195 21641 11204 21675
rect 11152 21632 11204 21641
rect 12440 21632 12492 21684
rect 19984 21675 20036 21684
rect 19984 21641 19993 21675
rect 19993 21641 20027 21675
rect 20027 21641 20036 21675
rect 19984 21632 20036 21641
rect 20720 21632 20772 21684
rect 21916 21632 21968 21684
rect 22376 21632 22428 21684
rect 23848 21632 23900 21684
rect 24492 21632 24544 21684
rect 25504 21675 25556 21684
rect 25504 21641 25513 21675
rect 25513 21641 25547 21675
rect 25547 21641 25556 21675
rect 25504 21632 25556 21641
rect 11704 21564 11756 21616
rect 1676 21539 1728 21548
rect 1676 21505 1685 21539
rect 1685 21505 1719 21539
rect 1719 21505 1728 21539
rect 1676 21496 1728 21505
rect 4160 21496 4212 21548
rect 4804 21539 4856 21548
rect 4804 21505 4813 21539
rect 4813 21505 4847 21539
rect 4847 21505 4856 21539
rect 4804 21496 4856 21505
rect 4988 21539 5040 21548
rect 4988 21505 4997 21539
rect 4997 21505 5031 21539
rect 5031 21505 5040 21539
rect 4988 21496 5040 21505
rect 10140 21496 10192 21548
rect 11244 21496 11296 21548
rect 1400 21471 1452 21480
rect 1400 21437 1409 21471
rect 1409 21437 1443 21471
rect 1443 21437 1452 21471
rect 1400 21428 1452 21437
rect 3056 21428 3108 21480
rect 3884 21471 3936 21480
rect 3884 21437 3893 21471
rect 3893 21437 3927 21471
rect 3927 21437 3936 21471
rect 3884 21428 3936 21437
rect 4068 21471 4120 21480
rect 4068 21437 4077 21471
rect 4077 21437 4111 21471
rect 4111 21437 4120 21471
rect 4068 21428 4120 21437
rect 8024 21471 8076 21480
rect 8024 21437 8033 21471
rect 8033 21437 8067 21471
rect 8067 21437 8076 21471
rect 8024 21428 8076 21437
rect 8668 21471 8720 21480
rect 2596 21292 2648 21344
rect 3976 21335 4028 21344
rect 3976 21301 3985 21335
rect 3985 21301 4019 21335
rect 4019 21301 4028 21335
rect 3976 21292 4028 21301
rect 5724 21292 5776 21344
rect 8208 21292 8260 21344
rect 8668 21437 8677 21471
rect 8677 21437 8711 21471
rect 8711 21437 8720 21471
rect 8668 21428 8720 21437
rect 8760 21428 8812 21480
rect 9404 21471 9456 21480
rect 9404 21437 9413 21471
rect 9413 21437 9447 21471
rect 9447 21437 9456 21471
rect 9404 21428 9456 21437
rect 10784 21428 10836 21480
rect 11796 21428 11848 21480
rect 12532 21564 12584 21616
rect 24768 21607 24820 21616
rect 9680 21403 9732 21412
rect 9680 21369 9689 21403
rect 9689 21369 9723 21403
rect 9723 21369 9732 21403
rect 9680 21360 9732 21369
rect 12532 21428 12584 21480
rect 24768 21573 24777 21607
rect 24777 21573 24811 21607
rect 24811 21573 24820 21607
rect 24768 21564 24820 21573
rect 14372 21539 14424 21548
rect 14372 21505 14381 21539
rect 14381 21505 14415 21539
rect 14415 21505 14424 21539
rect 14372 21496 14424 21505
rect 12900 21428 12952 21480
rect 13820 21471 13872 21480
rect 13820 21437 13829 21471
rect 13829 21437 13863 21471
rect 13863 21437 13872 21471
rect 13820 21428 13872 21437
rect 14740 21496 14792 21548
rect 19708 21496 19760 21548
rect 15016 21471 15068 21480
rect 9864 21292 9916 21344
rect 12440 21292 12492 21344
rect 14004 21360 14056 21412
rect 15016 21437 15025 21471
rect 15025 21437 15059 21471
rect 15059 21437 15068 21471
rect 15016 21428 15068 21437
rect 12808 21292 12860 21344
rect 17684 21428 17736 21480
rect 21824 21496 21876 21548
rect 21916 21496 21968 21548
rect 22652 21496 22704 21548
rect 29460 21632 29512 21684
rect 27252 21564 27304 21616
rect 22928 21471 22980 21480
rect 18696 21360 18748 21412
rect 22928 21437 22937 21471
rect 22937 21437 22971 21471
rect 22971 21437 22980 21471
rect 22928 21428 22980 21437
rect 23572 21428 23624 21480
rect 22468 21360 22520 21412
rect 23112 21360 23164 21412
rect 27068 21496 27120 21548
rect 24860 21471 24912 21480
rect 24860 21437 24869 21471
rect 24869 21437 24903 21471
rect 24903 21437 24912 21471
rect 24860 21428 24912 21437
rect 27988 21471 28040 21480
rect 27988 21437 27997 21471
rect 27997 21437 28031 21471
rect 28031 21437 28040 21471
rect 27988 21428 28040 21437
rect 28172 21428 28224 21480
rect 31208 21496 31260 21548
rect 31392 21496 31444 21548
rect 31852 21496 31904 21548
rect 32956 21496 33008 21548
rect 33600 21471 33652 21480
rect 33600 21437 33609 21471
rect 33609 21437 33643 21471
rect 33643 21437 33652 21471
rect 33600 21428 33652 21437
rect 25320 21360 25372 21412
rect 26424 21360 26476 21412
rect 32220 21360 32272 21412
rect 18512 21292 18564 21344
rect 22928 21292 22980 21344
rect 23940 21292 23992 21344
rect 26148 21292 26200 21344
rect 29000 21292 29052 21344
rect 32128 21335 32180 21344
rect 32128 21301 32137 21335
rect 32137 21301 32171 21335
rect 32171 21301 32180 21335
rect 32128 21292 32180 21301
rect 33416 21335 33468 21344
rect 33416 21301 33425 21335
rect 33425 21301 33459 21335
rect 33459 21301 33468 21335
rect 33416 21292 33468 21301
rect 12052 21190 12104 21242
rect 12116 21190 12168 21242
rect 12180 21190 12232 21242
rect 12244 21190 12296 21242
rect 23123 21190 23175 21242
rect 23187 21190 23239 21242
rect 23251 21190 23303 21242
rect 23315 21190 23367 21242
rect 4344 21088 4396 21140
rect 3976 21020 4028 21072
rect 3148 20995 3200 21004
rect 3148 20961 3157 20995
rect 3157 20961 3191 20995
rect 3191 20961 3200 20995
rect 3148 20952 3200 20961
rect 3332 20952 3384 21004
rect 6920 21088 6972 21140
rect 7288 21131 7340 21140
rect 7288 21097 7297 21131
rect 7297 21097 7331 21131
rect 7331 21097 7340 21131
rect 7288 21088 7340 21097
rect 8668 21088 8720 21140
rect 11428 21131 11480 21140
rect 5448 20952 5500 21004
rect 5540 20952 5592 21004
rect 8208 21063 8260 21072
rect 8208 21029 8217 21063
rect 8217 21029 8251 21063
rect 8251 21029 8260 21063
rect 8208 21020 8260 21029
rect 9312 21020 9364 21072
rect 9588 21020 9640 21072
rect 9864 21020 9916 21072
rect 6368 20995 6420 21004
rect 6368 20961 6377 20995
rect 6377 20961 6411 20995
rect 6411 20961 6420 20995
rect 6368 20952 6420 20961
rect 7012 20952 7064 21004
rect 11428 21097 11437 21131
rect 11437 21097 11471 21131
rect 11471 21097 11480 21131
rect 11428 21088 11480 21097
rect 11888 21088 11940 21140
rect 15016 21088 15068 21140
rect 17408 21088 17460 21140
rect 17684 21131 17736 21140
rect 17684 21097 17693 21131
rect 17693 21097 17727 21131
rect 17727 21097 17736 21131
rect 17684 21088 17736 21097
rect 4436 20884 4488 20936
rect 4528 20884 4580 20936
rect 2964 20859 3016 20868
rect 2964 20825 2973 20859
rect 2973 20825 3007 20859
rect 3007 20825 3016 20859
rect 2964 20816 3016 20825
rect 4620 20816 4672 20868
rect 8208 20884 8260 20936
rect 9588 20884 9640 20936
rect 9772 20884 9824 20936
rect 10968 20952 11020 21004
rect 11888 20995 11940 21004
rect 3976 20748 4028 20800
rect 6368 20748 6420 20800
rect 8392 20748 8444 20800
rect 10508 20748 10560 20800
rect 11888 20961 11897 20995
rect 11897 20961 11931 20995
rect 11931 20961 11940 20995
rect 11888 20952 11940 20961
rect 12808 21020 12860 21072
rect 33416 21088 33468 21140
rect 22468 21063 22520 21072
rect 12532 20952 12584 21004
rect 14556 20952 14608 21004
rect 15108 20952 15160 21004
rect 22468 21029 22477 21063
rect 22477 21029 22511 21063
rect 22511 21029 22520 21063
rect 22468 21020 22520 21029
rect 24032 21063 24084 21072
rect 24032 21029 24041 21063
rect 24041 21029 24075 21063
rect 24075 21029 24084 21063
rect 24032 21020 24084 21029
rect 24860 21020 24912 21072
rect 27436 21020 27488 21072
rect 32128 21063 32180 21072
rect 32128 21029 32137 21063
rect 32137 21029 32171 21063
rect 32171 21029 32180 21063
rect 32128 21020 32180 21029
rect 32588 21020 32640 21072
rect 16580 20995 16632 21004
rect 16580 20961 16614 20995
rect 16614 20961 16632 20995
rect 18696 20995 18748 21004
rect 16580 20952 16632 20961
rect 18696 20961 18705 20995
rect 18705 20961 18739 20995
rect 18739 20961 18748 20995
rect 18696 20952 18748 20961
rect 20352 20995 20404 21004
rect 20352 20961 20361 20995
rect 20361 20961 20395 20995
rect 20395 20961 20404 20995
rect 20352 20952 20404 20961
rect 22376 20995 22428 21004
rect 22376 20961 22385 20995
rect 22385 20961 22419 20995
rect 22419 20961 22428 20995
rect 22376 20952 22428 20961
rect 22744 20952 22796 21004
rect 12256 20884 12308 20936
rect 12440 20927 12492 20936
rect 12440 20893 12449 20927
rect 12449 20893 12483 20927
rect 12483 20893 12492 20927
rect 12440 20884 12492 20893
rect 14924 20927 14976 20936
rect 14924 20893 14933 20927
rect 14933 20893 14967 20927
rect 14967 20893 14976 20927
rect 14924 20884 14976 20893
rect 16304 20927 16356 20936
rect 16304 20893 16313 20927
rect 16313 20893 16347 20927
rect 16347 20893 16356 20927
rect 16304 20884 16356 20893
rect 19432 20884 19484 20936
rect 20996 20884 21048 20936
rect 23756 20952 23808 21004
rect 23940 20995 23992 21004
rect 23940 20961 23949 20995
rect 23949 20961 23983 20995
rect 23983 20961 23992 20995
rect 23940 20952 23992 20961
rect 25504 20952 25556 21004
rect 26148 20952 26200 21004
rect 26516 20995 26568 21004
rect 26516 20961 26525 20995
rect 26525 20961 26559 20995
rect 26559 20961 26568 20995
rect 26516 20952 26568 20961
rect 27252 20995 27304 21004
rect 27252 20961 27261 20995
rect 27261 20961 27295 20995
rect 27295 20961 27304 20995
rect 27252 20952 27304 20961
rect 29092 20995 29144 21004
rect 29092 20961 29110 20995
rect 29110 20961 29144 20995
rect 29092 20952 29144 20961
rect 30840 20995 30892 21004
rect 30840 20961 30849 20995
rect 30849 20961 30883 20995
rect 30883 20961 30892 20995
rect 30840 20952 30892 20961
rect 25228 20884 25280 20936
rect 25320 20884 25372 20936
rect 26424 20884 26476 20936
rect 19064 20816 19116 20868
rect 29368 20927 29420 20936
rect 29368 20893 29377 20927
rect 29377 20893 29411 20927
rect 29411 20893 29420 20927
rect 29368 20884 29420 20893
rect 29828 20884 29880 20936
rect 31208 20884 31260 20936
rect 31760 20884 31812 20936
rect 32220 20884 32272 20936
rect 12900 20748 12952 20800
rect 18328 20748 18380 20800
rect 18972 20748 19024 20800
rect 20168 20791 20220 20800
rect 20168 20757 20177 20791
rect 20177 20757 20211 20791
rect 20211 20757 20220 20791
rect 20168 20748 20220 20757
rect 23940 20748 23992 20800
rect 26608 20748 26660 20800
rect 27620 20748 27672 20800
rect 30472 20791 30524 20800
rect 30472 20757 30481 20791
rect 30481 20757 30515 20791
rect 30515 20757 30524 20791
rect 30472 20748 30524 20757
rect 6517 20646 6569 20698
rect 6581 20646 6633 20698
rect 6645 20646 6697 20698
rect 6709 20646 6761 20698
rect 17588 20646 17640 20698
rect 17652 20646 17704 20698
rect 17716 20646 17768 20698
rect 17780 20646 17832 20698
rect 28658 20646 28710 20698
rect 28722 20646 28774 20698
rect 28786 20646 28838 20698
rect 28850 20646 28902 20698
rect 3148 20544 3200 20596
rect 3332 20587 3384 20596
rect 3332 20553 3341 20587
rect 3341 20553 3375 20587
rect 3375 20553 3384 20587
rect 3332 20544 3384 20553
rect 4068 20544 4120 20596
rect 6920 20587 6972 20596
rect 6920 20553 6929 20587
rect 6929 20553 6963 20587
rect 6963 20553 6972 20587
rect 6920 20544 6972 20553
rect 8208 20544 8260 20596
rect 9680 20544 9732 20596
rect 11888 20544 11940 20596
rect 12348 20544 12400 20596
rect 19432 20587 19484 20596
rect 19432 20553 19441 20587
rect 19441 20553 19475 20587
rect 19475 20553 19484 20587
rect 19432 20544 19484 20553
rect 20168 20544 20220 20596
rect 23848 20544 23900 20596
rect 24768 20544 24820 20596
rect 25964 20587 26016 20596
rect 25964 20553 25973 20587
rect 25973 20553 26007 20587
rect 26007 20553 26016 20587
rect 25964 20544 26016 20553
rect 26056 20544 26108 20596
rect 29092 20544 29144 20596
rect 30840 20544 30892 20596
rect 1768 20451 1820 20460
rect 1768 20417 1777 20451
rect 1777 20417 1811 20451
rect 1811 20417 1820 20451
rect 1768 20408 1820 20417
rect 3976 20408 4028 20460
rect 8392 20451 8444 20460
rect 8392 20417 8401 20451
rect 8401 20417 8435 20451
rect 8435 20417 8444 20451
rect 8392 20408 8444 20417
rect 9404 20408 9456 20460
rect 3884 20383 3936 20392
rect 1952 20315 2004 20324
rect 1952 20281 1961 20315
rect 1961 20281 1995 20315
rect 1995 20281 2004 20315
rect 1952 20272 2004 20281
rect 3884 20349 3893 20383
rect 3893 20349 3927 20383
rect 3927 20349 3936 20383
rect 3884 20340 3936 20349
rect 4804 20340 4856 20392
rect 5448 20340 5500 20392
rect 5724 20383 5776 20392
rect 5724 20349 5733 20383
rect 5733 20349 5767 20383
rect 5767 20349 5776 20383
rect 5724 20340 5776 20349
rect 9956 20340 10008 20392
rect 10508 20383 10560 20392
rect 7012 20272 7064 20324
rect 8944 20272 8996 20324
rect 5080 20204 5132 20256
rect 10508 20349 10517 20383
rect 10517 20349 10551 20383
rect 10551 20349 10560 20383
rect 10508 20340 10560 20349
rect 13452 20476 13504 20528
rect 13544 20476 13596 20528
rect 11060 20383 11112 20392
rect 11060 20349 11069 20383
rect 11069 20349 11103 20383
rect 11103 20349 11112 20383
rect 11060 20340 11112 20349
rect 11336 20340 11388 20392
rect 12532 20340 12584 20392
rect 13176 20340 13228 20392
rect 13636 20340 13688 20392
rect 14004 20383 14056 20392
rect 14004 20349 14013 20383
rect 14013 20349 14047 20383
rect 14047 20349 14056 20383
rect 14004 20340 14056 20349
rect 10968 20272 11020 20324
rect 12440 20272 12492 20324
rect 13268 20272 13320 20324
rect 15844 20315 15896 20324
rect 15844 20281 15853 20315
rect 15853 20281 15887 20315
rect 15887 20281 15896 20315
rect 15844 20272 15896 20281
rect 16304 20408 16356 20460
rect 17316 20383 17368 20392
rect 17316 20349 17325 20383
rect 17325 20349 17359 20383
rect 17359 20349 17368 20383
rect 17316 20340 17368 20349
rect 17408 20340 17460 20392
rect 18328 20383 18380 20392
rect 18328 20349 18362 20383
rect 18362 20349 18380 20383
rect 18328 20340 18380 20349
rect 20996 20340 21048 20392
rect 27252 20476 27304 20528
rect 22192 20408 22244 20460
rect 22560 20408 22612 20460
rect 23020 20383 23072 20392
rect 23020 20349 23029 20383
rect 23029 20349 23063 20383
rect 23063 20349 23072 20383
rect 23020 20340 23072 20349
rect 23480 20383 23532 20392
rect 23480 20349 23489 20383
rect 23489 20349 23523 20383
rect 23523 20349 23532 20383
rect 23480 20340 23532 20349
rect 23756 20383 23808 20392
rect 23756 20349 23765 20383
rect 23765 20349 23799 20383
rect 23799 20349 23808 20383
rect 23756 20340 23808 20349
rect 23940 20408 23992 20460
rect 28264 20408 28316 20460
rect 29000 20408 29052 20460
rect 30472 20408 30524 20460
rect 16120 20272 16172 20324
rect 16764 20272 16816 20324
rect 22836 20315 22888 20324
rect 22836 20281 22845 20315
rect 22845 20281 22879 20315
rect 22879 20281 22888 20315
rect 22836 20272 22888 20281
rect 24032 20272 24084 20324
rect 25320 20340 25372 20392
rect 25780 20383 25832 20392
rect 25780 20349 25789 20383
rect 25789 20349 25823 20383
rect 25823 20349 25832 20383
rect 25780 20340 25832 20349
rect 26424 20383 26476 20392
rect 26424 20349 26433 20383
rect 26433 20349 26467 20383
rect 26467 20349 26476 20383
rect 26424 20340 26476 20349
rect 26608 20340 26660 20392
rect 28448 20383 28500 20392
rect 28448 20349 28457 20383
rect 28457 20349 28491 20383
rect 28491 20349 28500 20383
rect 28448 20340 28500 20349
rect 32036 20544 32088 20596
rect 32220 20340 32272 20392
rect 12992 20204 13044 20256
rect 13912 20204 13964 20256
rect 14096 20247 14148 20256
rect 14096 20213 14105 20247
rect 14105 20213 14139 20247
rect 14139 20213 14148 20247
rect 14096 20204 14148 20213
rect 14832 20204 14884 20256
rect 18420 20204 18472 20256
rect 19064 20204 19116 20256
rect 20168 20247 20220 20256
rect 20168 20213 20177 20247
rect 20177 20213 20211 20247
rect 20211 20213 20220 20247
rect 20168 20204 20220 20213
rect 23572 20204 23624 20256
rect 29828 20272 29880 20324
rect 32588 20272 32640 20324
rect 25596 20204 25648 20256
rect 27620 20204 27672 20256
rect 12052 20102 12104 20154
rect 12116 20102 12168 20154
rect 12180 20102 12232 20154
rect 12244 20102 12296 20154
rect 23123 20102 23175 20154
rect 23187 20102 23239 20154
rect 23251 20102 23303 20154
rect 23315 20102 23367 20154
rect 3056 20000 3108 20052
rect 3332 20000 3384 20052
rect 4160 20000 4212 20052
rect 5448 20000 5500 20052
rect 6828 20043 6880 20052
rect 2688 19864 2740 19916
rect 3332 19907 3384 19916
rect 2228 19839 2280 19848
rect 2228 19805 2237 19839
rect 2237 19805 2271 19839
rect 2271 19805 2280 19839
rect 2228 19796 2280 19805
rect 3332 19873 3341 19907
rect 3341 19873 3375 19907
rect 3375 19873 3384 19907
rect 3332 19864 3384 19873
rect 3884 19864 3936 19916
rect 5264 19932 5316 19984
rect 6828 20009 6837 20043
rect 6837 20009 6871 20043
rect 6871 20009 6880 20043
rect 6828 20000 6880 20009
rect 5080 19864 5132 19916
rect 5632 19864 5684 19916
rect 9680 19932 9732 19984
rect 15200 20000 15252 20052
rect 16580 20000 16632 20052
rect 9772 19907 9824 19916
rect 9772 19873 9781 19907
rect 9781 19873 9815 19907
rect 9815 19873 9824 19907
rect 9772 19864 9824 19873
rect 10140 19907 10192 19916
rect 10140 19873 10149 19907
rect 10149 19873 10183 19907
rect 10183 19873 10192 19907
rect 10140 19864 10192 19873
rect 12532 19975 12584 19984
rect 12532 19941 12541 19975
rect 12541 19941 12575 19975
rect 12575 19941 12584 19975
rect 12532 19932 12584 19941
rect 16304 19932 16356 19984
rect 19064 20000 19116 20052
rect 20352 20000 20404 20052
rect 10692 19907 10744 19916
rect 10692 19873 10701 19907
rect 10701 19873 10735 19907
rect 10735 19873 10744 19907
rect 10692 19864 10744 19873
rect 12256 19864 12308 19916
rect 12808 19864 12860 19916
rect 4712 19796 4764 19848
rect 7104 19796 7156 19848
rect 11796 19796 11848 19848
rect 14096 19864 14148 19916
rect 1952 19728 2004 19780
rect 1676 19660 1728 19712
rect 3148 19660 3200 19712
rect 4068 19660 4120 19712
rect 12900 19728 12952 19780
rect 15016 19907 15068 19916
rect 15016 19873 15025 19907
rect 15025 19873 15059 19907
rect 15059 19873 15068 19907
rect 15016 19864 15068 19873
rect 16764 19907 16816 19916
rect 16764 19873 16773 19907
rect 16773 19873 16807 19907
rect 16807 19873 16816 19907
rect 16764 19864 16816 19873
rect 18972 19932 19024 19984
rect 21364 19932 21416 19984
rect 25320 19932 25372 19984
rect 26516 20043 26568 20052
rect 26516 20009 26525 20043
rect 26525 20009 26559 20043
rect 26559 20009 26568 20043
rect 26516 20000 26568 20009
rect 14832 19660 14884 19712
rect 14924 19660 14976 19712
rect 16120 19728 16172 19780
rect 17316 19864 17368 19916
rect 17868 19907 17920 19916
rect 17868 19873 17877 19907
rect 17877 19873 17911 19907
rect 17911 19873 17920 19907
rect 17868 19864 17920 19873
rect 20260 19796 20312 19848
rect 20720 19796 20772 19848
rect 23020 19864 23072 19916
rect 24308 19907 24360 19916
rect 24308 19873 24317 19907
rect 24317 19873 24351 19907
rect 24351 19873 24360 19907
rect 24308 19864 24360 19873
rect 24768 19864 24820 19916
rect 25780 19864 25832 19916
rect 27620 19932 27672 19984
rect 32588 19932 32640 19984
rect 26424 19907 26476 19916
rect 26424 19873 26433 19907
rect 26433 19873 26467 19907
rect 26467 19873 26476 19907
rect 26424 19864 26476 19873
rect 27252 19907 27304 19916
rect 27252 19873 27261 19907
rect 27261 19873 27295 19907
rect 27295 19873 27304 19907
rect 27252 19864 27304 19873
rect 27344 19864 27396 19916
rect 18696 19728 18748 19780
rect 21640 19728 21692 19780
rect 25688 19796 25740 19848
rect 28264 19839 28316 19848
rect 28264 19805 28273 19839
rect 28273 19805 28307 19839
rect 28307 19805 28316 19839
rect 28264 19796 28316 19805
rect 28448 19839 28500 19848
rect 28448 19805 28457 19839
rect 28457 19805 28491 19839
rect 28491 19805 28500 19839
rect 28448 19796 28500 19805
rect 31760 19796 31812 19848
rect 32128 19839 32180 19848
rect 32128 19805 32137 19839
rect 32137 19805 32171 19839
rect 32171 19805 32180 19839
rect 32128 19796 32180 19805
rect 15752 19660 15804 19712
rect 16028 19660 16080 19712
rect 16580 19660 16632 19712
rect 22100 19703 22152 19712
rect 22100 19669 22109 19703
rect 22109 19669 22143 19703
rect 22143 19669 22152 19703
rect 22100 19660 22152 19669
rect 22652 19660 22704 19712
rect 29552 19660 29604 19712
rect 33600 19703 33652 19712
rect 33600 19669 33609 19703
rect 33609 19669 33643 19703
rect 33643 19669 33652 19703
rect 33600 19660 33652 19669
rect 6517 19558 6569 19610
rect 6581 19558 6633 19610
rect 6645 19558 6697 19610
rect 6709 19558 6761 19610
rect 17588 19558 17640 19610
rect 17652 19558 17704 19610
rect 17716 19558 17768 19610
rect 17780 19558 17832 19610
rect 28658 19558 28710 19610
rect 28722 19558 28774 19610
rect 28786 19558 28838 19610
rect 28850 19558 28902 19610
rect 3332 19456 3384 19508
rect 3976 19499 4028 19508
rect 3976 19465 3985 19499
rect 3985 19465 4019 19499
rect 4019 19465 4028 19499
rect 3976 19456 4028 19465
rect 4436 19456 4488 19508
rect 10508 19456 10560 19508
rect 12256 19499 12308 19508
rect 10692 19388 10744 19440
rect 12256 19465 12265 19499
rect 12265 19465 12299 19499
rect 12299 19465 12308 19499
rect 12256 19456 12308 19465
rect 13176 19499 13228 19508
rect 13176 19465 13185 19499
rect 13185 19465 13219 19499
rect 13219 19465 13228 19499
rect 13176 19456 13228 19465
rect 13544 19499 13596 19508
rect 13544 19465 13553 19499
rect 13553 19465 13587 19499
rect 13587 19465 13596 19499
rect 13544 19456 13596 19465
rect 14832 19456 14884 19508
rect 15844 19456 15896 19508
rect 21640 19456 21692 19508
rect 24308 19456 24360 19508
rect 27252 19456 27304 19508
rect 13820 19388 13872 19440
rect 14648 19388 14700 19440
rect 16028 19388 16080 19440
rect 32220 19388 32272 19440
rect 1676 19363 1728 19372
rect 1676 19329 1685 19363
rect 1685 19329 1719 19363
rect 1719 19329 1728 19363
rect 1676 19320 1728 19329
rect 5632 19363 5684 19372
rect 5632 19329 5641 19363
rect 5641 19329 5675 19363
rect 5675 19329 5684 19363
rect 5632 19320 5684 19329
rect 7104 19363 7156 19372
rect 7104 19329 7113 19363
rect 7113 19329 7147 19363
rect 7147 19329 7156 19363
rect 7104 19320 7156 19329
rect 1400 19295 1452 19304
rect 1400 19261 1409 19295
rect 1409 19261 1443 19295
rect 1443 19261 1452 19295
rect 1400 19252 1452 19261
rect 4528 19295 4580 19304
rect 2412 19184 2464 19236
rect 4528 19261 4537 19295
rect 4537 19261 4571 19295
rect 4571 19261 4580 19295
rect 4528 19252 4580 19261
rect 4712 19295 4764 19304
rect 4712 19261 4721 19295
rect 4721 19261 4755 19295
rect 4755 19261 4764 19295
rect 4712 19252 4764 19261
rect 5080 19252 5132 19304
rect 5540 19295 5592 19304
rect 5540 19261 5549 19295
rect 5549 19261 5583 19295
rect 5583 19261 5592 19295
rect 5540 19252 5592 19261
rect 4160 19116 4212 19168
rect 8944 19252 8996 19304
rect 9312 19252 9364 19304
rect 9588 19295 9640 19304
rect 9588 19261 9597 19295
rect 9597 19261 9631 19295
rect 9631 19261 9640 19295
rect 9588 19252 9640 19261
rect 10048 19295 10100 19304
rect 7012 19184 7064 19236
rect 8392 19116 8444 19168
rect 8484 19116 8536 19168
rect 10048 19261 10057 19295
rect 10057 19261 10091 19295
rect 10091 19261 10100 19295
rect 10048 19252 10100 19261
rect 9864 19184 9916 19236
rect 11796 19252 11848 19304
rect 11520 19184 11572 19236
rect 12900 19320 12952 19372
rect 13636 19320 13688 19372
rect 13360 19295 13412 19304
rect 10692 19116 10744 19168
rect 13360 19261 13369 19295
rect 13369 19261 13403 19295
rect 13403 19261 13412 19295
rect 13360 19252 13412 19261
rect 13452 19252 13504 19304
rect 13912 19252 13964 19304
rect 15752 19320 15804 19372
rect 20628 19320 20680 19372
rect 15476 19295 15528 19304
rect 15476 19261 15485 19295
rect 15485 19261 15519 19295
rect 15519 19261 15528 19295
rect 15476 19252 15528 19261
rect 15844 19295 15896 19304
rect 15844 19261 15853 19295
rect 15853 19261 15887 19295
rect 15887 19261 15896 19295
rect 15844 19252 15896 19261
rect 16120 19295 16172 19304
rect 16120 19261 16129 19295
rect 16129 19261 16163 19295
rect 16163 19261 16172 19295
rect 16120 19252 16172 19261
rect 19892 19295 19944 19304
rect 14004 19184 14056 19236
rect 15016 19184 15068 19236
rect 15292 19227 15344 19236
rect 15292 19193 15301 19227
rect 15301 19193 15335 19227
rect 15335 19193 15344 19227
rect 15292 19184 15344 19193
rect 14832 19116 14884 19168
rect 15108 19116 15160 19168
rect 15752 19184 15804 19236
rect 19892 19261 19901 19295
rect 19901 19261 19935 19295
rect 19935 19261 19944 19295
rect 19892 19252 19944 19261
rect 20352 19252 20404 19304
rect 20812 19294 20864 19346
rect 20904 19363 20956 19372
rect 20904 19329 20913 19363
rect 20913 19329 20947 19363
rect 20947 19329 20956 19363
rect 20904 19320 20956 19329
rect 22468 19320 22520 19372
rect 23572 19363 23624 19372
rect 23572 19329 23581 19363
rect 23581 19329 23615 19363
rect 23615 19329 23624 19363
rect 23572 19320 23624 19329
rect 30840 19320 30892 19372
rect 31208 19363 31260 19372
rect 31208 19329 31217 19363
rect 31217 19329 31251 19363
rect 31251 19329 31260 19363
rect 31208 19320 31260 19329
rect 33600 19320 33652 19372
rect 16580 19184 16632 19236
rect 17776 19184 17828 19236
rect 20720 19227 20772 19236
rect 20720 19193 20729 19227
rect 20729 19193 20763 19227
rect 20763 19193 20772 19227
rect 20720 19184 20772 19193
rect 20996 19295 21048 19304
rect 20996 19261 21005 19295
rect 21005 19261 21039 19295
rect 21039 19261 21048 19295
rect 20996 19252 21048 19261
rect 22100 19252 22152 19304
rect 22652 19295 22704 19304
rect 22652 19261 22661 19295
rect 22661 19261 22695 19295
rect 22695 19261 22704 19295
rect 22652 19252 22704 19261
rect 22744 19252 22796 19304
rect 25320 19252 25372 19304
rect 22560 19184 22612 19236
rect 23020 19184 23072 19236
rect 23664 19184 23716 19236
rect 25136 19184 25188 19236
rect 26608 19295 26660 19304
rect 26608 19261 26617 19295
rect 26617 19261 26651 19295
rect 26651 19261 26660 19295
rect 26608 19252 26660 19261
rect 27344 19252 27396 19304
rect 29552 19295 29604 19304
rect 29552 19261 29570 19295
rect 29570 19261 29604 19295
rect 29828 19295 29880 19304
rect 29552 19252 29604 19261
rect 29828 19261 29837 19295
rect 29837 19261 29871 19295
rect 29871 19261 29880 19295
rect 29828 19252 29880 19261
rect 31760 19252 31812 19304
rect 26976 19184 27028 19236
rect 15936 19159 15988 19168
rect 15936 19125 15945 19159
rect 15945 19125 15979 19159
rect 15979 19125 15988 19159
rect 15936 19116 15988 19125
rect 19800 19116 19852 19168
rect 20444 19116 20496 19168
rect 25228 19116 25280 19168
rect 25688 19159 25740 19168
rect 25688 19125 25697 19159
rect 25697 19125 25731 19159
rect 25731 19125 25740 19159
rect 25688 19116 25740 19125
rect 26240 19116 26292 19168
rect 28448 19159 28500 19168
rect 28448 19125 28457 19159
rect 28457 19125 28491 19159
rect 28491 19125 28500 19159
rect 28448 19116 28500 19125
rect 30748 19116 30800 19168
rect 32220 19116 32272 19168
rect 33048 19159 33100 19168
rect 33048 19125 33057 19159
rect 33057 19125 33091 19159
rect 33091 19125 33100 19159
rect 33048 19116 33100 19125
rect 12052 19014 12104 19066
rect 12116 19014 12168 19066
rect 12180 19014 12232 19066
rect 12244 19014 12296 19066
rect 23123 19014 23175 19066
rect 23187 19014 23239 19066
rect 23251 19014 23303 19066
rect 23315 19014 23367 19066
rect 2228 18912 2280 18964
rect 4528 18912 4580 18964
rect 5540 18912 5592 18964
rect 9864 18912 9916 18964
rect 10048 18912 10100 18964
rect 2688 18844 2740 18896
rect 4160 18844 4212 18896
rect 5080 18887 5132 18896
rect 3332 18819 3384 18828
rect 3332 18785 3341 18819
rect 3341 18785 3375 18819
rect 3375 18785 3384 18819
rect 3332 18776 3384 18785
rect 5080 18853 5089 18887
rect 5089 18853 5123 18887
rect 5123 18853 5132 18887
rect 5080 18844 5132 18853
rect 10968 18844 11020 18896
rect 15476 18844 15528 18896
rect 5724 18819 5776 18828
rect 5724 18785 5733 18819
rect 5733 18785 5767 18819
rect 5767 18785 5776 18819
rect 5724 18776 5776 18785
rect 6184 18776 6236 18828
rect 6828 18776 6880 18828
rect 8484 18819 8536 18828
rect 8484 18785 8493 18819
rect 8493 18785 8527 18819
rect 8527 18785 8536 18819
rect 8484 18776 8536 18785
rect 9680 18819 9732 18828
rect 9680 18785 9689 18819
rect 9689 18785 9723 18819
rect 9723 18785 9732 18819
rect 9680 18776 9732 18785
rect 10692 18776 10744 18828
rect 11336 18776 11388 18828
rect 11520 18819 11572 18828
rect 11520 18785 11529 18819
rect 11529 18785 11563 18819
rect 11563 18785 11572 18819
rect 11520 18776 11572 18785
rect 10232 18708 10284 18760
rect 10600 18708 10652 18760
rect 11704 18708 11756 18760
rect 13360 18776 13412 18828
rect 13636 18819 13688 18828
rect 13636 18785 13645 18819
rect 13645 18785 13679 18819
rect 13679 18785 13688 18819
rect 13636 18776 13688 18785
rect 13912 18776 13964 18828
rect 12440 18751 12492 18760
rect 12440 18717 12449 18751
rect 12449 18717 12483 18751
rect 12483 18717 12492 18751
rect 12716 18751 12768 18760
rect 12440 18708 12492 18717
rect 12716 18717 12725 18751
rect 12725 18717 12759 18751
rect 12759 18717 12768 18751
rect 12716 18708 12768 18717
rect 13544 18708 13596 18760
rect 4068 18640 4120 18692
rect 10324 18640 10376 18692
rect 10416 18640 10468 18692
rect 14924 18776 14976 18828
rect 16304 18844 16356 18896
rect 17408 18912 17460 18964
rect 17776 18912 17828 18964
rect 18052 18844 18104 18896
rect 19892 18912 19944 18964
rect 25136 18912 25188 18964
rect 26516 18912 26568 18964
rect 32128 18912 32180 18964
rect 33600 18912 33652 18964
rect 15200 18751 15252 18760
rect 15200 18717 15209 18751
rect 15209 18717 15243 18751
rect 15243 18717 15252 18751
rect 15200 18708 15252 18717
rect 16028 18776 16080 18828
rect 19708 18776 19760 18828
rect 19892 18819 19944 18828
rect 19892 18785 19901 18819
rect 19901 18785 19935 18819
rect 19935 18785 19944 18819
rect 19892 18776 19944 18785
rect 20168 18819 20220 18828
rect 20168 18785 20177 18819
rect 20177 18785 20211 18819
rect 20211 18785 20220 18819
rect 20168 18776 20220 18785
rect 25320 18776 25372 18828
rect 26332 18844 26384 18896
rect 30748 18887 30800 18896
rect 30748 18853 30757 18887
rect 30757 18853 30791 18887
rect 30791 18853 30800 18887
rect 30748 18844 30800 18853
rect 32588 18844 32640 18896
rect 26148 18819 26200 18828
rect 26148 18785 26157 18819
rect 26157 18785 26191 18819
rect 26191 18785 26200 18819
rect 26148 18776 26200 18785
rect 26700 18819 26752 18828
rect 26700 18785 26709 18819
rect 26709 18785 26743 18819
rect 26743 18785 26752 18819
rect 26700 18776 26752 18785
rect 27252 18776 27304 18828
rect 28172 18819 28224 18828
rect 28172 18785 28181 18819
rect 28181 18785 28215 18819
rect 28215 18785 28224 18819
rect 28172 18776 28224 18785
rect 18972 18751 19024 18760
rect 18972 18717 18981 18751
rect 18981 18717 19015 18751
rect 19015 18717 19024 18751
rect 18972 18708 19024 18717
rect 19616 18751 19668 18760
rect 19616 18717 19625 18751
rect 19625 18717 19659 18751
rect 19659 18717 19668 18751
rect 19616 18708 19668 18717
rect 19800 18751 19852 18760
rect 19800 18717 19809 18751
rect 19809 18717 19843 18751
rect 19843 18717 19852 18751
rect 19800 18708 19852 18717
rect 20352 18751 20404 18760
rect 20352 18717 20361 18751
rect 20361 18717 20395 18751
rect 20395 18717 20404 18751
rect 20352 18708 20404 18717
rect 28448 18776 28500 18828
rect 29828 18776 29880 18828
rect 31208 18708 31260 18760
rect 32220 18751 32272 18760
rect 5724 18572 5776 18624
rect 16856 18640 16908 18692
rect 17868 18640 17920 18692
rect 10692 18615 10744 18624
rect 10692 18581 10701 18615
rect 10701 18581 10735 18615
rect 10735 18581 10744 18615
rect 10692 18572 10744 18581
rect 12808 18572 12860 18624
rect 17040 18572 17092 18624
rect 19524 18640 19576 18692
rect 25964 18640 26016 18692
rect 27896 18683 27948 18692
rect 27896 18649 27905 18683
rect 27905 18649 27939 18683
rect 27939 18649 27948 18683
rect 27896 18640 27948 18649
rect 32220 18717 32229 18751
rect 32229 18717 32263 18751
rect 32263 18717 32272 18751
rect 32220 18708 32272 18717
rect 19064 18572 19116 18624
rect 25412 18615 25464 18624
rect 25412 18581 25421 18615
rect 25421 18581 25455 18615
rect 25455 18581 25464 18615
rect 27160 18615 27212 18624
rect 25412 18572 25464 18581
rect 27160 18581 27169 18615
rect 27169 18581 27203 18615
rect 27203 18581 27212 18615
rect 27160 18572 27212 18581
rect 28080 18572 28132 18624
rect 6517 18470 6569 18522
rect 6581 18470 6633 18522
rect 6645 18470 6697 18522
rect 6709 18470 6761 18522
rect 17588 18470 17640 18522
rect 17652 18470 17704 18522
rect 17716 18470 17768 18522
rect 17780 18470 17832 18522
rect 28658 18470 28710 18522
rect 28722 18470 28774 18522
rect 28786 18470 28838 18522
rect 28850 18470 28902 18522
rect 8208 18368 8260 18420
rect 9588 18368 9640 18420
rect 10692 18368 10744 18420
rect 10968 18368 11020 18420
rect 12348 18368 12400 18420
rect 12440 18368 12492 18420
rect 12900 18368 12952 18420
rect 15016 18368 15068 18420
rect 15752 18368 15804 18420
rect 17408 18368 17460 18420
rect 2504 18207 2556 18216
rect 2504 18173 2513 18207
rect 2513 18173 2547 18207
rect 2547 18173 2556 18207
rect 2504 18164 2556 18173
rect 2780 18164 2832 18216
rect 3240 18164 3292 18216
rect 5080 18232 5132 18284
rect 3056 18139 3108 18148
rect 3056 18105 3065 18139
rect 3065 18105 3099 18139
rect 3099 18105 3108 18139
rect 3056 18096 3108 18105
rect 4252 18139 4304 18148
rect 4252 18105 4261 18139
rect 4261 18105 4295 18139
rect 4295 18105 4304 18139
rect 5264 18207 5316 18216
rect 5264 18173 5273 18207
rect 5273 18173 5307 18207
rect 5307 18173 5316 18207
rect 5264 18164 5316 18173
rect 6828 18164 6880 18216
rect 7288 18164 7340 18216
rect 12256 18300 12308 18352
rect 9864 18232 9916 18284
rect 4252 18096 4304 18105
rect 6184 18096 6236 18148
rect 3884 18071 3936 18080
rect 3884 18037 3893 18071
rect 3893 18037 3927 18071
rect 3927 18037 3936 18071
rect 3884 18028 3936 18037
rect 4160 18028 4212 18080
rect 4988 18028 5040 18080
rect 8484 18028 8536 18080
rect 9588 18207 9640 18216
rect 9588 18173 9597 18207
rect 9597 18173 9631 18207
rect 9631 18173 9640 18207
rect 9588 18164 9640 18173
rect 10048 18096 10100 18148
rect 9956 18028 10008 18080
rect 11152 18207 11204 18216
rect 11152 18173 11161 18207
rect 11161 18173 11195 18207
rect 11195 18173 11204 18207
rect 11152 18164 11204 18173
rect 11060 18071 11112 18080
rect 11060 18037 11069 18071
rect 11069 18037 11103 18071
rect 11103 18037 11112 18071
rect 11060 18028 11112 18037
rect 12716 18232 12768 18284
rect 14832 18275 14884 18284
rect 14832 18241 14841 18275
rect 14841 18241 14875 18275
rect 14875 18241 14884 18275
rect 14832 18232 14884 18241
rect 16672 18300 16724 18352
rect 19892 18368 19944 18420
rect 22652 18411 22704 18420
rect 19708 18300 19760 18352
rect 22652 18377 22661 18411
rect 22661 18377 22695 18411
rect 22695 18377 22704 18411
rect 22652 18368 22704 18377
rect 26148 18368 26200 18420
rect 27804 18411 27856 18420
rect 27804 18377 27813 18411
rect 27813 18377 27847 18411
rect 27847 18377 27856 18411
rect 27804 18368 27856 18377
rect 30564 18411 30616 18420
rect 30564 18377 30573 18411
rect 30573 18377 30607 18411
rect 30607 18377 30616 18411
rect 30564 18368 30616 18377
rect 31576 18368 31628 18420
rect 20260 18300 20312 18352
rect 12440 18207 12492 18216
rect 12440 18173 12449 18207
rect 12449 18173 12483 18207
rect 12483 18173 12492 18207
rect 12808 18207 12860 18216
rect 12440 18164 12492 18173
rect 12808 18173 12817 18207
rect 12817 18173 12851 18207
rect 12851 18173 12860 18207
rect 12808 18164 12860 18173
rect 13268 18207 13320 18216
rect 13268 18173 13277 18207
rect 13277 18173 13311 18207
rect 13311 18173 13320 18207
rect 13268 18164 13320 18173
rect 13728 18207 13780 18216
rect 13728 18173 13737 18207
rect 13737 18173 13771 18207
rect 13771 18173 13780 18207
rect 13728 18164 13780 18173
rect 15016 18207 15068 18216
rect 15016 18173 15025 18207
rect 15025 18173 15059 18207
rect 15059 18173 15068 18207
rect 15016 18164 15068 18173
rect 15476 18164 15528 18216
rect 18052 18232 18104 18284
rect 19064 18275 19116 18284
rect 19064 18241 19073 18275
rect 19073 18241 19107 18275
rect 19107 18241 19116 18275
rect 19064 18232 19116 18241
rect 22744 18232 22796 18284
rect 18604 18096 18656 18148
rect 21088 18096 21140 18148
rect 21364 18139 21416 18148
rect 21364 18105 21373 18139
rect 21373 18105 21407 18139
rect 21407 18105 21416 18139
rect 21364 18096 21416 18105
rect 23664 18096 23716 18148
rect 24124 18139 24176 18148
rect 24124 18105 24133 18139
rect 24133 18105 24167 18139
rect 24167 18105 24176 18139
rect 24124 18096 24176 18105
rect 27160 18232 27212 18284
rect 25412 18164 25464 18216
rect 27804 18164 27856 18216
rect 28080 18207 28132 18216
rect 28080 18173 28089 18207
rect 28089 18173 28123 18207
rect 28123 18173 28132 18207
rect 28080 18164 28132 18173
rect 30656 18164 30708 18216
rect 30932 18164 30984 18216
rect 29828 18096 29880 18148
rect 12716 18028 12768 18080
rect 15384 18028 15436 18080
rect 15844 18028 15896 18080
rect 18972 18028 19024 18080
rect 21272 18028 21324 18080
rect 12052 17926 12104 17978
rect 12116 17926 12168 17978
rect 12180 17926 12232 17978
rect 12244 17926 12296 17978
rect 23123 17926 23175 17978
rect 23187 17926 23239 17978
rect 23251 17926 23303 17978
rect 23315 17926 23367 17978
rect 2504 17824 2556 17876
rect 2872 17824 2924 17876
rect 8392 17824 8444 17876
rect 9680 17824 9732 17876
rect 3056 17799 3108 17808
rect 3056 17765 3065 17799
rect 3065 17765 3099 17799
rect 3099 17765 3108 17799
rect 3056 17756 3108 17765
rect 2596 17688 2648 17740
rect 4344 17731 4396 17740
rect 4344 17697 4353 17731
rect 4353 17697 4387 17731
rect 4387 17697 4396 17731
rect 4344 17688 4396 17697
rect 4712 17756 4764 17808
rect 5264 17756 5316 17808
rect 17224 17824 17276 17876
rect 21364 17824 21416 17876
rect 24124 17824 24176 17876
rect 27896 17824 27948 17876
rect 14924 17756 14976 17808
rect 2872 17663 2924 17672
rect 2872 17629 2881 17663
rect 2881 17629 2915 17663
rect 2915 17629 2924 17663
rect 2872 17620 2924 17629
rect 2596 17484 2648 17536
rect 4896 17484 4948 17536
rect 5908 17731 5960 17740
rect 5908 17697 5917 17731
rect 5917 17697 5951 17731
rect 5951 17697 5960 17731
rect 5908 17688 5960 17697
rect 6184 17731 6236 17740
rect 6184 17697 6193 17731
rect 6193 17697 6227 17731
rect 6227 17697 6236 17731
rect 6184 17688 6236 17697
rect 6368 17731 6420 17740
rect 6368 17697 6377 17731
rect 6377 17697 6411 17731
rect 6411 17697 6420 17731
rect 6368 17688 6420 17697
rect 7472 17731 7524 17740
rect 7472 17697 7481 17731
rect 7481 17697 7515 17731
rect 7515 17697 7524 17731
rect 7472 17688 7524 17697
rect 10416 17731 10468 17740
rect 10416 17697 10425 17731
rect 10425 17697 10459 17731
rect 10459 17697 10468 17731
rect 10416 17688 10468 17697
rect 11888 17688 11940 17740
rect 12992 17731 13044 17740
rect 12992 17697 13001 17731
rect 13001 17697 13035 17731
rect 13035 17697 13044 17731
rect 12992 17688 13044 17697
rect 14648 17688 14700 17740
rect 15384 17756 15436 17808
rect 15936 17756 15988 17808
rect 16120 17756 16172 17808
rect 15476 17688 15528 17740
rect 17408 17688 17460 17740
rect 20720 17688 20772 17740
rect 21272 17731 21324 17740
rect 21272 17697 21281 17731
rect 21281 17697 21315 17731
rect 21315 17697 21324 17731
rect 21272 17688 21324 17697
rect 22100 17756 22152 17808
rect 22652 17731 22704 17740
rect 10784 17620 10836 17672
rect 7196 17552 7248 17604
rect 11612 17552 11664 17604
rect 12716 17620 12768 17672
rect 13728 17620 13780 17672
rect 15200 17620 15252 17672
rect 22652 17697 22661 17731
rect 22661 17697 22695 17731
rect 22695 17697 22704 17731
rect 22652 17688 22704 17697
rect 22836 17731 22888 17740
rect 22836 17697 22845 17731
rect 22845 17697 22879 17731
rect 22879 17697 22888 17731
rect 22836 17688 22888 17697
rect 26792 17756 26844 17808
rect 27620 17756 27672 17808
rect 32588 17756 32640 17808
rect 27988 17731 28040 17740
rect 26424 17620 26476 17672
rect 27988 17697 27997 17731
rect 27997 17697 28031 17731
rect 28031 17697 28040 17731
rect 27988 17688 28040 17697
rect 31760 17688 31812 17740
rect 27804 17663 27856 17672
rect 27804 17629 27813 17663
rect 27813 17629 27847 17663
rect 27847 17629 27856 17663
rect 27804 17620 27856 17629
rect 28264 17663 28316 17672
rect 28264 17629 28273 17663
rect 28273 17629 28307 17663
rect 28307 17629 28316 17663
rect 28264 17620 28316 17629
rect 32128 17663 32180 17672
rect 32128 17629 32137 17663
rect 32137 17629 32171 17663
rect 32171 17629 32180 17663
rect 32128 17620 32180 17629
rect 7380 17527 7432 17536
rect 7380 17493 7389 17527
rect 7389 17493 7423 17527
rect 7423 17493 7432 17527
rect 7380 17484 7432 17493
rect 9588 17484 9640 17536
rect 11520 17484 11572 17536
rect 11796 17484 11848 17536
rect 12348 17484 12400 17536
rect 13084 17484 13136 17536
rect 13636 17484 13688 17536
rect 14832 17484 14884 17536
rect 17224 17484 17276 17536
rect 19616 17484 19668 17536
rect 19984 17484 20036 17536
rect 22744 17484 22796 17536
rect 33508 17484 33560 17536
rect 6517 17382 6569 17434
rect 6581 17382 6633 17434
rect 6645 17382 6697 17434
rect 6709 17382 6761 17434
rect 17588 17382 17640 17434
rect 17652 17382 17704 17434
rect 17716 17382 17768 17434
rect 17780 17382 17832 17434
rect 28658 17382 28710 17434
rect 28722 17382 28774 17434
rect 28786 17382 28838 17434
rect 28850 17382 28902 17434
rect 2780 17323 2832 17332
rect 2780 17289 2789 17323
rect 2789 17289 2823 17323
rect 2823 17289 2832 17323
rect 4712 17323 4764 17332
rect 2780 17280 2832 17289
rect 4712 17289 4721 17323
rect 4721 17289 4755 17323
rect 4755 17289 4764 17323
rect 4712 17280 4764 17289
rect 4896 17323 4948 17332
rect 4896 17289 4905 17323
rect 4905 17289 4939 17323
rect 4939 17289 4948 17323
rect 4896 17280 4948 17289
rect 5908 17280 5960 17332
rect 9956 17323 10008 17332
rect 7380 17187 7432 17196
rect 7380 17153 7389 17187
rect 7389 17153 7423 17187
rect 7423 17153 7432 17187
rect 7380 17144 7432 17153
rect 2596 17119 2648 17128
rect 2596 17085 2605 17119
rect 2605 17085 2639 17119
rect 2639 17085 2648 17119
rect 2596 17076 2648 17085
rect 4252 17076 4304 17128
rect 4804 17076 4856 17128
rect 5632 17119 5684 17128
rect 2872 17008 2924 17060
rect 5632 17085 5641 17119
rect 5641 17085 5675 17119
rect 5675 17085 5684 17119
rect 5632 17076 5684 17085
rect 7196 17119 7248 17128
rect 7196 17085 7205 17119
rect 7205 17085 7239 17119
rect 7239 17085 7248 17119
rect 9956 17289 9965 17323
rect 9965 17289 9999 17323
rect 9999 17289 10008 17323
rect 9956 17280 10008 17289
rect 11152 17323 11204 17332
rect 11152 17289 11161 17323
rect 11161 17289 11195 17323
rect 11195 17289 11204 17323
rect 11152 17280 11204 17289
rect 25136 17280 25188 17332
rect 28172 17280 28224 17332
rect 13728 17212 13780 17264
rect 8484 17187 8536 17196
rect 8484 17153 8493 17187
rect 8493 17153 8527 17187
rect 8527 17153 8536 17187
rect 8484 17144 8536 17153
rect 11704 17144 11756 17196
rect 7196 17076 7248 17085
rect 12532 17119 12584 17128
rect 6368 17008 6420 17060
rect 8392 17008 8444 17060
rect 6828 16983 6880 16992
rect 6828 16949 6837 16983
rect 6837 16949 6871 16983
rect 6871 16949 6880 16983
rect 6828 16940 6880 16949
rect 7288 16983 7340 16992
rect 7288 16949 7297 16983
rect 7297 16949 7331 16983
rect 7331 16949 7340 16983
rect 12532 17085 12541 17119
rect 12541 17085 12575 17119
rect 12575 17085 12584 17119
rect 12532 17076 12584 17085
rect 13084 17119 13136 17128
rect 13084 17085 13093 17119
rect 13093 17085 13127 17119
rect 13127 17085 13136 17119
rect 13084 17076 13136 17085
rect 15108 17187 15160 17196
rect 15108 17153 15117 17187
rect 15117 17153 15151 17187
rect 15151 17153 15160 17187
rect 15108 17144 15160 17153
rect 16120 17144 16172 17196
rect 17316 17144 17368 17196
rect 13636 17119 13688 17128
rect 13636 17085 13645 17119
rect 13645 17085 13679 17119
rect 13679 17085 13688 17119
rect 13636 17076 13688 17085
rect 12440 17051 12492 17060
rect 12440 17017 12449 17051
rect 12449 17017 12483 17051
rect 12483 17017 12492 17051
rect 12440 17008 12492 17017
rect 13544 17008 13596 17060
rect 15016 17119 15068 17128
rect 15016 17085 15025 17119
rect 15025 17085 15059 17119
rect 15059 17085 15068 17119
rect 15016 17076 15068 17085
rect 15384 17008 15436 17060
rect 15752 17051 15804 17060
rect 15752 17017 15761 17051
rect 15761 17017 15795 17051
rect 15795 17017 15804 17051
rect 15752 17008 15804 17017
rect 17224 17008 17276 17060
rect 7288 16940 7340 16949
rect 12808 16940 12860 16992
rect 13452 16940 13504 16992
rect 17132 16940 17184 16992
rect 24584 17144 24636 17196
rect 25596 17187 25648 17196
rect 25596 17153 25605 17187
rect 25605 17153 25639 17187
rect 25639 17153 25648 17187
rect 25596 17144 25648 17153
rect 18972 17051 19024 17060
rect 18972 17017 18981 17051
rect 18981 17017 19015 17051
rect 19015 17017 19024 17051
rect 18972 17008 19024 17017
rect 19984 17076 20036 17128
rect 22100 17076 22152 17128
rect 24952 17119 25004 17128
rect 24952 17085 24961 17119
rect 24961 17085 24995 17119
rect 24995 17085 25004 17119
rect 24952 17076 25004 17085
rect 26240 17076 26292 17128
rect 26700 17119 26752 17128
rect 20904 17008 20956 17060
rect 23664 17008 23716 17060
rect 25964 17051 26016 17060
rect 18604 16940 18656 16992
rect 19800 16983 19852 16992
rect 19800 16949 19809 16983
rect 19809 16949 19843 16983
rect 19843 16949 19852 16983
rect 19800 16940 19852 16949
rect 23756 16940 23808 16992
rect 24584 16940 24636 16992
rect 25964 17017 25973 17051
rect 25973 17017 26007 17051
rect 26007 17017 26016 17051
rect 25964 17008 26016 17017
rect 26700 17085 26709 17119
rect 26709 17085 26743 17119
rect 26743 17085 26752 17119
rect 26700 17076 26752 17085
rect 27988 17119 28040 17128
rect 27988 17085 27997 17119
rect 27997 17085 28031 17119
rect 28031 17085 28040 17119
rect 27988 17076 28040 17085
rect 28264 17076 28316 17128
rect 30288 17212 30340 17264
rect 32588 17212 32640 17264
rect 30564 17187 30616 17196
rect 30564 17153 30573 17187
rect 30573 17153 30607 17187
rect 30607 17153 30616 17187
rect 30564 17144 30616 17153
rect 31208 17119 31260 17128
rect 25688 16940 25740 16992
rect 26148 16940 26200 16992
rect 31208 17085 31217 17119
rect 31217 17085 31251 17119
rect 31251 17085 31260 17119
rect 31208 17076 31260 17085
rect 32036 17119 32088 17128
rect 29092 17051 29144 17060
rect 29092 17017 29101 17051
rect 29101 17017 29135 17051
rect 29135 17017 29144 17051
rect 29092 17008 29144 17017
rect 30840 17008 30892 17060
rect 32036 17085 32045 17119
rect 32045 17085 32079 17119
rect 32079 17085 32088 17119
rect 32036 17076 32088 17085
rect 33140 17076 33192 17128
rect 32220 17008 32272 17060
rect 33600 17051 33652 17060
rect 33600 17017 33609 17051
rect 33609 17017 33643 17051
rect 33643 17017 33652 17051
rect 33600 17008 33652 17017
rect 29000 16940 29052 16992
rect 31024 16983 31076 16992
rect 31024 16949 31033 16983
rect 31033 16949 31067 16983
rect 31067 16949 31076 16983
rect 31024 16940 31076 16949
rect 31944 16983 31996 16992
rect 31944 16949 31953 16983
rect 31953 16949 31987 16983
rect 31987 16949 31996 16983
rect 31944 16940 31996 16949
rect 12052 16838 12104 16890
rect 12116 16838 12168 16890
rect 12180 16838 12232 16890
rect 12244 16838 12296 16890
rect 23123 16838 23175 16890
rect 23187 16838 23239 16890
rect 23251 16838 23303 16890
rect 23315 16838 23367 16890
rect 4344 16736 4396 16788
rect 7288 16736 7340 16788
rect 11888 16779 11940 16788
rect 11888 16745 11897 16779
rect 11897 16745 11931 16779
rect 11931 16745 11940 16779
rect 11888 16736 11940 16745
rect 12532 16779 12584 16788
rect 12532 16745 12541 16779
rect 12541 16745 12575 16779
rect 12575 16745 12584 16779
rect 12532 16736 12584 16745
rect 15108 16736 15160 16788
rect 3424 16668 3476 16720
rect 6828 16711 6880 16720
rect 6828 16677 6862 16711
rect 6862 16677 6880 16711
rect 6828 16668 6880 16677
rect 2964 16643 3016 16652
rect 2964 16609 2968 16643
rect 2968 16609 3002 16643
rect 3002 16609 3016 16643
rect 2964 16600 3016 16609
rect 3332 16643 3384 16652
rect 3332 16609 3341 16643
rect 3341 16609 3375 16643
rect 3375 16609 3384 16643
rect 3332 16600 3384 16609
rect 4160 16600 4212 16652
rect 5632 16643 5684 16652
rect 5632 16609 5641 16643
rect 5641 16609 5675 16643
rect 5675 16609 5684 16643
rect 10048 16668 10100 16720
rect 5632 16600 5684 16609
rect 11520 16600 11572 16652
rect 12348 16600 12400 16652
rect 15016 16668 15068 16720
rect 12716 16600 12768 16652
rect 13268 16600 13320 16652
rect 13452 16643 13504 16652
rect 13452 16609 13461 16643
rect 13461 16609 13495 16643
rect 13495 16609 13504 16643
rect 13452 16600 13504 16609
rect 13912 16600 13964 16652
rect 14556 16600 14608 16652
rect 14832 16600 14884 16652
rect 17408 16736 17460 16788
rect 20996 16736 21048 16788
rect 17316 16668 17368 16720
rect 16396 16643 16448 16652
rect 6368 16532 6420 16584
rect 13544 16507 13596 16516
rect 13544 16473 13553 16507
rect 13553 16473 13587 16507
rect 13587 16473 13596 16507
rect 13544 16464 13596 16473
rect 16396 16609 16405 16643
rect 16405 16609 16439 16643
rect 16439 16609 16448 16643
rect 16396 16600 16448 16609
rect 17224 16643 17276 16652
rect 17224 16609 17233 16643
rect 17233 16609 17267 16643
rect 17267 16609 17276 16643
rect 17224 16600 17276 16609
rect 18604 16600 18656 16652
rect 15476 16464 15528 16516
rect 17316 16532 17368 16584
rect 20444 16600 20496 16652
rect 20628 16600 20680 16652
rect 22100 16600 22152 16652
rect 21088 16532 21140 16584
rect 21916 16532 21968 16584
rect 23664 16600 23716 16652
rect 25228 16643 25280 16652
rect 25228 16609 25237 16643
rect 25237 16609 25271 16643
rect 25271 16609 25280 16643
rect 25228 16600 25280 16609
rect 26516 16736 26568 16788
rect 32128 16736 32180 16788
rect 25688 16600 25740 16652
rect 26240 16600 26292 16652
rect 28540 16668 28592 16720
rect 30840 16711 30892 16720
rect 30840 16677 30849 16711
rect 30849 16677 30883 16711
rect 30883 16677 30892 16711
rect 30840 16668 30892 16677
rect 30564 16643 30616 16652
rect 26424 16532 26476 16584
rect 30564 16609 30573 16643
rect 30573 16609 30607 16643
rect 30607 16609 30616 16643
rect 30564 16600 30616 16609
rect 30748 16643 30800 16652
rect 30748 16609 30757 16643
rect 30757 16609 30791 16643
rect 30791 16609 30800 16643
rect 30748 16600 30800 16609
rect 31208 16600 31260 16652
rect 31392 16643 31444 16652
rect 31392 16609 31401 16643
rect 31401 16609 31435 16643
rect 31435 16609 31444 16643
rect 31392 16600 31444 16609
rect 31576 16643 31628 16652
rect 31576 16609 31585 16643
rect 31585 16609 31619 16643
rect 31619 16609 31628 16643
rect 31576 16600 31628 16609
rect 31944 16668 31996 16720
rect 32220 16668 32272 16720
rect 31852 16600 31904 16652
rect 32036 16532 32088 16584
rect 33508 16643 33560 16652
rect 33508 16609 33517 16643
rect 33517 16609 33551 16643
rect 33551 16609 33560 16643
rect 33508 16600 33560 16609
rect 20812 16464 20864 16516
rect 24768 16464 24820 16516
rect 26056 16464 26108 16516
rect 3056 16396 3108 16448
rect 15936 16396 15988 16448
rect 16948 16396 17000 16448
rect 19984 16396 20036 16448
rect 20444 16396 20496 16448
rect 26516 16396 26568 16448
rect 6517 16294 6569 16346
rect 6581 16294 6633 16346
rect 6645 16294 6697 16346
rect 6709 16294 6761 16346
rect 17588 16294 17640 16346
rect 17652 16294 17704 16346
rect 17716 16294 17768 16346
rect 17780 16294 17832 16346
rect 28658 16294 28710 16346
rect 28722 16294 28774 16346
rect 28786 16294 28838 16346
rect 28850 16294 28902 16346
rect 4804 16235 4856 16244
rect 4804 16201 4813 16235
rect 4813 16201 4847 16235
rect 4847 16201 4856 16235
rect 4804 16192 4856 16201
rect 14096 16235 14148 16244
rect 14096 16201 14105 16235
rect 14105 16201 14139 16235
rect 14139 16201 14148 16235
rect 14096 16192 14148 16201
rect 14648 16192 14700 16244
rect 16396 16192 16448 16244
rect 18972 16192 19024 16244
rect 19524 16235 19576 16244
rect 19524 16201 19533 16235
rect 19533 16201 19567 16235
rect 19567 16201 19576 16235
rect 19524 16192 19576 16201
rect 20628 16192 20680 16244
rect 20904 16192 20956 16244
rect 11336 16124 11388 16176
rect 3424 16099 3476 16108
rect 3424 16065 3433 16099
rect 3433 16065 3467 16099
rect 3467 16065 3476 16099
rect 3424 16056 3476 16065
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 4160 16031 4212 16040
rect 4160 15997 4169 16031
rect 4169 15997 4203 16031
rect 4203 15997 4212 16031
rect 4160 15988 4212 15997
rect 10140 16056 10192 16108
rect 5172 16031 5224 16040
rect 5172 15997 5181 16031
rect 5181 15997 5215 16031
rect 5215 15997 5224 16031
rect 5172 15988 5224 15997
rect 6368 15988 6420 16040
rect 6644 15988 6696 16040
rect 10876 16031 10928 16040
rect 10876 15997 10885 16031
rect 10885 15997 10919 16031
rect 10919 15997 10928 16031
rect 10876 15988 10928 15997
rect 12900 16124 12952 16176
rect 16948 16124 17000 16176
rect 19984 16124 20036 16176
rect 13636 16056 13688 16108
rect 14832 16056 14884 16108
rect 13360 15988 13412 16040
rect 15936 15988 15988 16040
rect 17132 16056 17184 16108
rect 19800 16056 19852 16108
rect 20996 16099 21048 16108
rect 20996 16065 21005 16099
rect 21005 16065 21039 16099
rect 21039 16065 21048 16099
rect 20996 16056 21048 16065
rect 22468 16192 22520 16244
rect 26240 16235 26292 16244
rect 26240 16201 26249 16235
rect 26249 16201 26283 16235
rect 26283 16201 26292 16235
rect 26240 16192 26292 16201
rect 21732 16056 21784 16108
rect 25228 16056 25280 16108
rect 28264 16192 28316 16244
rect 29092 16192 29144 16244
rect 1676 15963 1728 15972
rect 1676 15929 1685 15963
rect 1685 15929 1719 15963
rect 1719 15929 1728 15963
rect 1676 15920 1728 15929
rect 2688 15920 2740 15972
rect 7564 15963 7616 15972
rect 7564 15929 7573 15963
rect 7573 15929 7607 15963
rect 7607 15929 7616 15963
rect 7564 15920 7616 15929
rect 8024 15920 8076 15972
rect 8852 15920 8904 15972
rect 8208 15852 8260 15904
rect 10876 15852 10928 15904
rect 12440 15852 12492 15904
rect 12900 15852 12952 15904
rect 13176 15852 13228 15904
rect 13728 15852 13780 15904
rect 13912 15852 13964 15904
rect 15752 15920 15804 15972
rect 17316 15920 17368 15972
rect 19524 15920 19576 15972
rect 15568 15852 15620 15904
rect 16212 15852 16264 15904
rect 20536 15920 20588 15972
rect 20720 15920 20772 15972
rect 23020 15988 23072 16040
rect 23480 16031 23532 16040
rect 23480 15997 23489 16031
rect 23489 15997 23523 16031
rect 23523 15997 23532 16031
rect 23480 15988 23532 15997
rect 25596 15988 25648 16040
rect 26332 16031 26384 16040
rect 22744 15920 22796 15972
rect 25320 15963 25372 15972
rect 25320 15929 25329 15963
rect 25329 15929 25363 15963
rect 25363 15929 25372 15963
rect 25320 15920 25372 15929
rect 26332 15997 26341 16031
rect 26341 15997 26375 16031
rect 26375 15997 26384 16031
rect 26332 15988 26384 15997
rect 28540 15988 28592 16040
rect 29184 15988 29236 16040
rect 31024 16124 31076 16176
rect 31576 16056 31628 16108
rect 30656 15988 30708 16040
rect 31392 15988 31444 16040
rect 31852 15988 31904 16040
rect 33600 16031 33652 16040
rect 33600 15997 33609 16031
rect 33609 15997 33643 16031
rect 33643 15997 33652 16031
rect 33600 15988 33652 15997
rect 30840 15920 30892 15972
rect 31208 15920 31260 15972
rect 20812 15852 20864 15904
rect 22008 15852 22060 15904
rect 32128 15895 32180 15904
rect 32128 15861 32137 15895
rect 32137 15861 32171 15895
rect 32171 15861 32180 15895
rect 32128 15852 32180 15861
rect 12052 15750 12104 15802
rect 12116 15750 12168 15802
rect 12180 15750 12232 15802
rect 12244 15750 12296 15802
rect 23123 15750 23175 15802
rect 23187 15750 23239 15802
rect 23251 15750 23303 15802
rect 23315 15750 23367 15802
rect 1676 15648 1728 15700
rect 2688 15580 2740 15632
rect 7012 15648 7064 15700
rect 8024 15648 8076 15700
rect 9772 15648 9824 15700
rect 7288 15580 7340 15632
rect 7472 15580 7524 15632
rect 9680 15623 9732 15632
rect 9680 15589 9689 15623
rect 9689 15589 9723 15623
rect 9723 15589 9732 15623
rect 9680 15580 9732 15589
rect 15384 15648 15436 15700
rect 10968 15580 11020 15632
rect 3056 15555 3108 15564
rect 3056 15521 3065 15555
rect 3065 15521 3099 15555
rect 3099 15521 3108 15555
rect 3056 15512 3108 15521
rect 3424 15512 3476 15564
rect 8208 15512 8260 15564
rect 10876 15512 10928 15564
rect 2964 15444 3016 15496
rect 4068 15444 4120 15496
rect 6368 15487 6420 15496
rect 6368 15453 6377 15487
rect 6377 15453 6411 15487
rect 6411 15453 6420 15487
rect 6368 15444 6420 15453
rect 6644 15487 6696 15496
rect 6644 15453 6653 15487
rect 6653 15453 6687 15487
rect 6687 15453 6696 15487
rect 6644 15444 6696 15453
rect 7840 15487 7892 15496
rect 7840 15453 7849 15487
rect 7849 15453 7883 15487
rect 7883 15453 7892 15487
rect 7840 15444 7892 15453
rect 4528 15308 4580 15360
rect 5172 15308 5224 15360
rect 6000 15308 6052 15360
rect 8300 15419 8352 15428
rect 8300 15385 8309 15419
rect 8309 15385 8343 15419
rect 8343 15385 8352 15419
rect 8300 15376 8352 15385
rect 11244 15512 11296 15564
rect 11336 15487 11388 15496
rect 11336 15453 11345 15487
rect 11345 15453 11379 15487
rect 11379 15453 11388 15487
rect 11336 15444 11388 15453
rect 13084 15580 13136 15632
rect 17316 15623 17368 15632
rect 17316 15589 17325 15623
rect 17325 15589 17359 15623
rect 17359 15589 17368 15623
rect 17316 15580 17368 15589
rect 12900 15512 12952 15564
rect 13360 15512 13412 15564
rect 13728 15512 13780 15564
rect 15568 15555 15620 15564
rect 15568 15521 15577 15555
rect 15577 15521 15611 15555
rect 15611 15521 15620 15555
rect 15568 15512 15620 15521
rect 16580 15512 16632 15564
rect 17224 15555 17276 15564
rect 17224 15521 17233 15555
rect 17233 15521 17267 15555
rect 17267 15521 17276 15555
rect 17224 15512 17276 15521
rect 20536 15648 20588 15700
rect 20720 15648 20772 15700
rect 21916 15648 21968 15700
rect 23480 15691 23532 15700
rect 22008 15623 22060 15632
rect 22008 15589 22017 15623
rect 22017 15589 22051 15623
rect 22051 15589 22060 15623
rect 22008 15580 22060 15589
rect 23480 15657 23489 15691
rect 23489 15657 23523 15691
rect 23523 15657 23532 15691
rect 23480 15648 23532 15657
rect 30840 15648 30892 15700
rect 17868 15512 17920 15564
rect 21732 15555 21784 15564
rect 21732 15521 21741 15555
rect 21741 15521 21775 15555
rect 21775 15521 21784 15555
rect 21732 15512 21784 15521
rect 25872 15580 25924 15632
rect 26056 15580 26108 15632
rect 25688 15512 25740 15564
rect 27988 15580 28040 15632
rect 26608 15512 26660 15564
rect 13452 15444 13504 15496
rect 16672 15444 16724 15496
rect 19064 15444 19116 15496
rect 25228 15487 25280 15496
rect 25228 15453 25237 15487
rect 25237 15453 25271 15487
rect 25271 15453 25280 15487
rect 25228 15444 25280 15453
rect 26332 15444 26384 15496
rect 27712 15512 27764 15564
rect 32036 15648 32088 15700
rect 33600 15691 33652 15700
rect 33600 15657 33609 15691
rect 33609 15657 33643 15691
rect 33643 15657 33652 15691
rect 33600 15648 33652 15657
rect 31852 15580 31904 15632
rect 32588 15580 32640 15632
rect 27620 15487 27672 15496
rect 12808 15376 12860 15428
rect 7472 15351 7524 15360
rect 7472 15317 7481 15351
rect 7481 15317 7515 15351
rect 7515 15317 7524 15351
rect 7472 15308 7524 15317
rect 10508 15308 10560 15360
rect 11796 15308 11848 15360
rect 12716 15308 12768 15360
rect 15752 15351 15804 15360
rect 15752 15317 15761 15351
rect 15761 15317 15795 15351
rect 15795 15317 15804 15351
rect 15752 15308 15804 15317
rect 17408 15308 17460 15360
rect 23940 15308 23992 15360
rect 25320 15351 25372 15360
rect 25320 15317 25329 15351
rect 25329 15317 25363 15351
rect 25363 15317 25372 15351
rect 25320 15308 25372 15317
rect 26056 15351 26108 15360
rect 26056 15317 26065 15351
rect 26065 15317 26099 15351
rect 26099 15317 26108 15351
rect 26056 15308 26108 15317
rect 26792 15308 26844 15360
rect 27620 15453 27629 15487
rect 27629 15453 27663 15487
rect 27663 15453 27672 15487
rect 27620 15444 27672 15453
rect 31760 15444 31812 15496
rect 31024 15351 31076 15360
rect 31024 15317 31033 15351
rect 31033 15317 31067 15351
rect 31067 15317 31076 15351
rect 31024 15308 31076 15317
rect 31208 15351 31260 15360
rect 31208 15317 31217 15351
rect 31217 15317 31251 15351
rect 31251 15317 31260 15351
rect 31208 15308 31260 15317
rect 6517 15206 6569 15258
rect 6581 15206 6633 15258
rect 6645 15206 6697 15258
rect 6709 15206 6761 15258
rect 17588 15206 17640 15258
rect 17652 15206 17704 15258
rect 17716 15206 17768 15258
rect 17780 15206 17832 15258
rect 28658 15206 28710 15258
rect 28722 15206 28774 15258
rect 28786 15206 28838 15258
rect 28850 15206 28902 15258
rect 10048 15104 10100 15156
rect 3424 15036 3476 15088
rect 4068 15011 4120 15020
rect 4068 14977 4077 15011
rect 4077 14977 4111 15011
rect 4111 14977 4120 15011
rect 11060 15036 11112 15088
rect 17408 15104 17460 15156
rect 17960 15104 18012 15156
rect 21824 15104 21876 15156
rect 4068 14968 4120 14977
rect 5080 14968 5132 15020
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 10784 15011 10836 15020
rect 10784 14977 10793 15011
rect 10793 14977 10827 15011
rect 10827 14977 10836 15011
rect 10784 14968 10836 14977
rect 13636 14968 13688 15020
rect 16396 14968 16448 15020
rect 22468 15036 22520 15088
rect 22284 14968 22336 15020
rect 24952 15104 25004 15156
rect 25780 15104 25832 15156
rect 25872 15104 25924 15156
rect 27712 15104 27764 15156
rect 30748 15147 30800 15156
rect 30748 15113 30757 15147
rect 30757 15113 30791 15147
rect 30791 15113 30800 15147
rect 30748 15104 30800 15113
rect 31852 15147 31904 15156
rect 31852 15113 31861 15147
rect 31861 15113 31895 15147
rect 31895 15113 31904 15147
rect 31852 15104 31904 15113
rect 26792 15011 26844 15020
rect 26792 14977 26801 15011
rect 26801 14977 26835 15011
rect 26835 14977 26844 15011
rect 26792 14968 26844 14977
rect 27620 14968 27672 15020
rect 29000 15011 29052 15020
rect 29000 14977 29009 15011
rect 29009 14977 29043 15011
rect 29043 14977 29052 15011
rect 29000 14968 29052 14977
rect 31668 14968 31720 15020
rect 1400 14943 1452 14952
rect 1400 14909 1409 14943
rect 1409 14909 1443 14943
rect 1443 14909 1452 14943
rect 1400 14900 1452 14909
rect 3332 14900 3384 14952
rect 4252 14900 4304 14952
rect 5172 14900 5224 14952
rect 7840 14943 7892 14952
rect 2688 14832 2740 14884
rect 4160 14832 4212 14884
rect 4528 14832 4580 14884
rect 7840 14909 7849 14943
rect 7849 14909 7883 14943
rect 7883 14909 7892 14943
rect 7840 14900 7892 14909
rect 8208 14943 8260 14952
rect 8208 14909 8217 14943
rect 8217 14909 8251 14943
rect 8251 14909 8260 14943
rect 8208 14900 8260 14909
rect 11888 14900 11940 14952
rect 13084 14943 13136 14952
rect 13084 14909 13093 14943
rect 13093 14909 13127 14943
rect 13127 14909 13136 14943
rect 13084 14900 13136 14909
rect 13452 14943 13504 14952
rect 13452 14909 13461 14943
rect 13461 14909 13495 14943
rect 13495 14909 13504 14943
rect 13452 14900 13504 14909
rect 15476 14943 15528 14952
rect 9772 14832 9824 14884
rect 15476 14909 15485 14943
rect 15485 14909 15519 14943
rect 15519 14909 15528 14943
rect 15476 14900 15528 14909
rect 16212 14900 16264 14952
rect 17316 14943 17368 14952
rect 17316 14909 17325 14943
rect 17325 14909 17359 14943
rect 17359 14909 17368 14943
rect 17316 14900 17368 14909
rect 20444 14900 20496 14952
rect 21732 14900 21784 14952
rect 25320 14900 25372 14952
rect 26516 14943 26568 14952
rect 26516 14909 26525 14943
rect 26525 14909 26559 14943
rect 26559 14909 26568 14943
rect 26516 14900 26568 14909
rect 30932 14900 30984 14952
rect 31392 14943 31444 14952
rect 31392 14909 31401 14943
rect 31401 14909 31435 14943
rect 31435 14909 31444 14943
rect 31392 14900 31444 14909
rect 31576 14900 31628 14952
rect 32128 14943 32180 14952
rect 32128 14909 32137 14943
rect 32137 14909 32171 14943
rect 32171 14909 32180 14943
rect 32128 14900 32180 14909
rect 15660 14832 15712 14884
rect 16672 14832 16724 14884
rect 20720 14832 20772 14884
rect 29276 14875 29328 14884
rect 29276 14841 29285 14875
rect 29285 14841 29319 14875
rect 29319 14841 29328 14875
rect 29276 14832 29328 14841
rect 30288 14832 30340 14884
rect 31760 14832 31812 14884
rect 5448 14764 5500 14816
rect 7288 14807 7340 14816
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 11244 14764 11296 14816
rect 17408 14764 17460 14816
rect 19064 14807 19116 14816
rect 19064 14773 19073 14807
rect 19073 14773 19107 14807
rect 19107 14773 19116 14807
rect 19064 14764 19116 14773
rect 20260 14764 20312 14816
rect 21456 14807 21508 14816
rect 21456 14773 21465 14807
rect 21465 14773 21499 14807
rect 21499 14773 21508 14807
rect 21456 14764 21508 14773
rect 32220 14764 32272 14816
rect 12052 14662 12104 14714
rect 12116 14662 12168 14714
rect 12180 14662 12232 14714
rect 12244 14662 12296 14714
rect 23123 14662 23175 14714
rect 23187 14662 23239 14714
rect 23251 14662 23303 14714
rect 23315 14662 23367 14714
rect 3424 14560 3476 14612
rect 4068 14560 4120 14612
rect 5172 14603 5224 14612
rect 5172 14569 5181 14603
rect 5181 14569 5215 14603
rect 5215 14569 5224 14603
rect 5172 14560 5224 14569
rect 4160 14492 4212 14544
rect 4528 14492 4580 14544
rect 7288 14560 7340 14612
rect 7564 14560 7616 14612
rect 12716 14560 12768 14612
rect 16580 14560 16632 14612
rect 5448 14492 5500 14544
rect 5080 14467 5132 14476
rect 5080 14433 5089 14467
rect 5089 14433 5123 14467
rect 5123 14433 5132 14467
rect 8300 14492 8352 14544
rect 12808 14492 12860 14544
rect 5080 14424 5132 14433
rect 7472 14467 7524 14476
rect 7472 14433 7481 14467
rect 7481 14433 7515 14467
rect 7515 14433 7524 14467
rect 7472 14424 7524 14433
rect 3332 14331 3384 14340
rect 3332 14297 3341 14331
rect 3341 14297 3375 14331
rect 3375 14297 3384 14331
rect 3332 14288 3384 14297
rect 4160 14288 4212 14340
rect 6368 14288 6420 14340
rect 11520 14424 11572 14476
rect 12256 14424 12308 14476
rect 12624 14424 12676 14476
rect 13452 14492 13504 14544
rect 15292 14424 15344 14476
rect 15752 14424 15804 14476
rect 18420 14492 18472 14544
rect 20904 14560 20956 14612
rect 21732 14603 21784 14612
rect 21732 14569 21741 14603
rect 21741 14569 21775 14603
rect 21775 14569 21784 14603
rect 22284 14603 22336 14612
rect 21732 14560 21784 14569
rect 20260 14535 20312 14544
rect 20260 14501 20269 14535
rect 20269 14501 20303 14535
rect 20303 14501 20312 14535
rect 20260 14492 20312 14501
rect 20720 14492 20772 14544
rect 16764 14467 16816 14476
rect 16764 14433 16773 14467
rect 16773 14433 16807 14467
rect 16807 14433 16816 14467
rect 16764 14424 16816 14433
rect 17960 14424 18012 14476
rect 18696 14424 18748 14476
rect 18788 14467 18840 14476
rect 18788 14433 18797 14467
rect 18797 14433 18831 14467
rect 18831 14433 18840 14467
rect 18788 14424 18840 14433
rect 18972 14467 19024 14476
rect 18972 14433 18981 14467
rect 18981 14433 19015 14467
rect 19015 14433 19024 14467
rect 19984 14467 20036 14476
rect 18972 14424 19024 14433
rect 19984 14433 19993 14467
rect 19993 14433 20027 14467
rect 20027 14433 20036 14467
rect 19984 14424 20036 14433
rect 22284 14569 22293 14603
rect 22293 14569 22327 14603
rect 22327 14569 22336 14603
rect 22284 14560 22336 14569
rect 25228 14560 25280 14612
rect 23020 14535 23072 14544
rect 22284 14424 22336 14476
rect 23020 14501 23029 14535
rect 23029 14501 23063 14535
rect 23063 14501 23072 14535
rect 23020 14492 23072 14501
rect 24400 14424 24452 14476
rect 26608 14560 26660 14612
rect 27988 14560 28040 14612
rect 29276 14560 29328 14612
rect 25780 14424 25832 14476
rect 26148 14492 26200 14544
rect 32036 14492 32088 14544
rect 30748 14467 30800 14476
rect 11612 14356 11664 14408
rect 13084 14356 13136 14408
rect 15476 14399 15528 14408
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 18236 14356 18288 14408
rect 30748 14433 30757 14467
rect 30757 14433 30791 14467
rect 30791 14433 30800 14467
rect 30748 14424 30800 14433
rect 31944 14424 31996 14476
rect 32220 14467 32272 14476
rect 32220 14433 32229 14467
rect 32229 14433 32263 14467
rect 32263 14433 32272 14467
rect 32220 14424 32272 14433
rect 33232 14424 33284 14476
rect 16856 14288 16908 14340
rect 19064 14288 19116 14340
rect 26608 14356 26660 14408
rect 23204 14331 23256 14340
rect 23204 14297 23213 14331
rect 23213 14297 23247 14331
rect 23247 14297 23256 14331
rect 23204 14288 23256 14297
rect 25872 14288 25924 14340
rect 12716 14220 12768 14272
rect 13544 14263 13596 14272
rect 13544 14229 13553 14263
rect 13553 14229 13587 14263
rect 13587 14229 13596 14263
rect 13544 14220 13596 14229
rect 15016 14263 15068 14272
rect 15016 14229 15025 14263
rect 15025 14229 15059 14263
rect 15059 14229 15068 14263
rect 15016 14220 15068 14229
rect 18236 14263 18288 14272
rect 18236 14229 18245 14263
rect 18245 14229 18279 14263
rect 18279 14229 18288 14263
rect 23756 14263 23808 14272
rect 18236 14220 18288 14229
rect 23756 14229 23765 14263
rect 23765 14229 23799 14263
rect 23799 14229 23808 14263
rect 23756 14220 23808 14229
rect 24952 14220 25004 14272
rect 27620 14220 27672 14272
rect 33324 14220 33376 14272
rect 6517 14118 6569 14170
rect 6581 14118 6633 14170
rect 6645 14118 6697 14170
rect 6709 14118 6761 14170
rect 17588 14118 17640 14170
rect 17652 14118 17704 14170
rect 17716 14118 17768 14170
rect 17780 14118 17832 14170
rect 28658 14118 28710 14170
rect 28722 14118 28774 14170
rect 28786 14118 28838 14170
rect 28850 14118 28902 14170
rect 13176 14016 13228 14068
rect 13636 14016 13688 14068
rect 15292 14059 15344 14068
rect 15292 14025 15301 14059
rect 15301 14025 15335 14059
rect 15335 14025 15344 14059
rect 15292 14016 15344 14025
rect 15660 14016 15712 14068
rect 17316 14016 17368 14068
rect 12900 13880 12952 13932
rect 5448 13855 5500 13864
rect 5448 13821 5457 13855
rect 5457 13821 5491 13855
rect 5491 13821 5500 13855
rect 5448 13812 5500 13821
rect 6000 13812 6052 13864
rect 7840 13812 7892 13864
rect 7932 13812 7984 13864
rect 11612 13812 11664 13864
rect 12256 13855 12308 13864
rect 12256 13821 12265 13855
rect 12265 13821 12299 13855
rect 12299 13821 12308 13855
rect 12256 13812 12308 13821
rect 12992 13855 13044 13864
rect 12992 13821 13001 13855
rect 13001 13821 13035 13855
rect 13035 13821 13044 13855
rect 12992 13812 13044 13821
rect 13544 13812 13596 13864
rect 15384 13812 15436 13864
rect 17408 13948 17460 14000
rect 19984 14016 20036 14068
rect 18972 13948 19024 14000
rect 21824 14016 21876 14068
rect 25596 14016 25648 14068
rect 26608 14059 26660 14068
rect 26608 14025 26617 14059
rect 26617 14025 26651 14059
rect 26651 14025 26660 14059
rect 26608 14016 26660 14025
rect 22468 13948 22520 14000
rect 15752 13812 15804 13864
rect 16212 13855 16264 13864
rect 16212 13821 16221 13855
rect 16221 13821 16255 13855
rect 16255 13821 16264 13855
rect 16212 13812 16264 13821
rect 16396 13855 16448 13864
rect 16396 13821 16405 13855
rect 16405 13821 16439 13855
rect 16439 13821 16448 13855
rect 16396 13812 16448 13821
rect 18236 13855 18288 13864
rect 18236 13821 18270 13855
rect 18270 13821 18288 13855
rect 18236 13812 18288 13821
rect 20812 13812 20864 13864
rect 22284 13880 22336 13932
rect 24400 13923 24452 13932
rect 24400 13889 24409 13923
rect 24409 13889 24443 13923
rect 24443 13889 24452 13923
rect 24400 13880 24452 13889
rect 21732 13812 21784 13864
rect 20904 13744 20956 13796
rect 26516 13855 26568 13864
rect 26516 13821 26525 13855
rect 26525 13821 26559 13855
rect 26559 13821 26568 13855
rect 26516 13812 26568 13821
rect 27988 13812 28040 13864
rect 31944 13855 31996 13864
rect 22928 13787 22980 13796
rect 22928 13753 22937 13787
rect 22937 13753 22971 13787
rect 22971 13753 22980 13787
rect 22928 13744 22980 13753
rect 23204 13744 23256 13796
rect 4068 13676 4120 13728
rect 4988 13676 5040 13728
rect 5356 13676 5408 13728
rect 6920 13719 6972 13728
rect 6920 13685 6929 13719
rect 6929 13685 6963 13719
rect 6963 13685 6972 13719
rect 6920 13676 6972 13685
rect 8760 13719 8812 13728
rect 8760 13685 8769 13719
rect 8769 13685 8803 13719
rect 8803 13685 8812 13719
rect 8760 13676 8812 13685
rect 9128 13719 9180 13728
rect 9128 13685 9137 13719
rect 9137 13685 9171 13719
rect 9171 13685 9180 13719
rect 9128 13676 9180 13685
rect 9588 13676 9640 13728
rect 12900 13676 12952 13728
rect 13912 13676 13964 13728
rect 15384 13676 15436 13728
rect 16120 13676 16172 13728
rect 20996 13719 21048 13728
rect 20996 13685 21005 13719
rect 21005 13685 21039 13719
rect 21039 13685 21048 13719
rect 20996 13676 21048 13685
rect 22836 13676 22888 13728
rect 25044 13744 25096 13796
rect 28540 13744 28592 13796
rect 30932 13787 30984 13796
rect 30932 13753 30941 13787
rect 30941 13753 30975 13787
rect 30975 13753 30984 13787
rect 30932 13744 30984 13753
rect 25964 13676 26016 13728
rect 29460 13719 29512 13728
rect 29460 13685 29469 13719
rect 29469 13685 29503 13719
rect 29503 13685 29512 13719
rect 29460 13676 29512 13685
rect 31944 13821 31953 13855
rect 31953 13821 31987 13855
rect 31987 13821 31996 13855
rect 31944 13812 31996 13821
rect 32220 13812 32272 13864
rect 33232 13855 33284 13864
rect 33232 13821 33241 13855
rect 33241 13821 33275 13855
rect 33275 13821 33284 13855
rect 33232 13812 33284 13821
rect 31760 13787 31812 13796
rect 31760 13753 31769 13787
rect 31769 13753 31803 13787
rect 31803 13753 31812 13787
rect 31760 13744 31812 13753
rect 31852 13676 31904 13728
rect 33416 13719 33468 13728
rect 33416 13685 33425 13719
rect 33425 13685 33459 13719
rect 33459 13685 33468 13719
rect 33416 13676 33468 13685
rect 12052 13574 12104 13626
rect 12116 13574 12168 13626
rect 12180 13574 12232 13626
rect 12244 13574 12296 13626
rect 23123 13574 23175 13626
rect 23187 13574 23239 13626
rect 23251 13574 23303 13626
rect 23315 13574 23367 13626
rect 7840 13472 7892 13524
rect 7012 13404 7064 13456
rect 12716 13515 12768 13524
rect 12716 13481 12725 13515
rect 12725 13481 12759 13515
rect 12759 13481 12768 13515
rect 12716 13472 12768 13481
rect 12808 13515 12860 13524
rect 12808 13481 12817 13515
rect 12817 13481 12851 13515
rect 12851 13481 12860 13515
rect 12808 13472 12860 13481
rect 2872 13379 2924 13388
rect 2872 13345 2881 13379
rect 2881 13345 2915 13379
rect 2915 13345 2924 13379
rect 2872 13336 2924 13345
rect 8668 13336 8720 13388
rect 2964 13311 3016 13320
rect 2964 13277 2973 13311
rect 2973 13277 3007 13311
rect 3007 13277 3016 13311
rect 2964 13268 3016 13277
rect 3056 13268 3108 13320
rect 4712 13268 4764 13320
rect 6000 13311 6052 13320
rect 6000 13277 6009 13311
rect 6009 13277 6043 13311
rect 6043 13277 6052 13311
rect 6000 13268 6052 13277
rect 6920 13268 6972 13320
rect 7012 13268 7064 13320
rect 8024 13268 8076 13320
rect 9956 13268 10008 13320
rect 10784 13268 10836 13320
rect 10968 13268 11020 13320
rect 11612 13336 11664 13388
rect 8852 13200 8904 13252
rect 12900 13311 12952 13320
rect 12900 13277 12909 13311
rect 12909 13277 12943 13311
rect 12943 13277 12952 13311
rect 12900 13268 12952 13277
rect 13544 13404 13596 13456
rect 13636 13336 13688 13388
rect 15200 13472 15252 13524
rect 20720 13472 20772 13524
rect 15016 13447 15068 13456
rect 15016 13413 15025 13447
rect 15025 13413 15059 13447
rect 15059 13413 15068 13447
rect 15016 13404 15068 13413
rect 15292 13404 15344 13456
rect 16764 13404 16816 13456
rect 22928 13472 22980 13524
rect 28540 13472 28592 13524
rect 26976 13447 27028 13456
rect 26976 13413 26985 13447
rect 26985 13413 27019 13447
rect 27019 13413 27028 13447
rect 26976 13404 27028 13413
rect 30380 13404 30432 13456
rect 32220 13472 32272 13524
rect 32588 13404 32640 13456
rect 16304 13336 16356 13388
rect 17408 13336 17460 13388
rect 18236 13379 18288 13388
rect 18236 13345 18245 13379
rect 18245 13345 18279 13379
rect 18279 13345 18288 13379
rect 18236 13336 18288 13345
rect 18420 13379 18472 13388
rect 18420 13345 18429 13379
rect 18429 13345 18463 13379
rect 18463 13345 18472 13379
rect 18420 13336 18472 13345
rect 18696 13336 18748 13388
rect 18972 13336 19024 13388
rect 22744 13379 22796 13388
rect 22744 13345 22753 13379
rect 22753 13345 22787 13379
rect 22787 13345 22796 13379
rect 22744 13336 22796 13345
rect 22836 13379 22888 13388
rect 22836 13345 22845 13379
rect 22845 13345 22879 13379
rect 22879 13345 22888 13379
rect 22836 13336 22888 13345
rect 26148 13336 26200 13388
rect 28172 13336 28224 13388
rect 29552 13336 29604 13388
rect 31024 13336 31076 13388
rect 15384 13268 15436 13320
rect 15476 13268 15528 13320
rect 16028 13268 16080 13320
rect 1768 13132 1820 13184
rect 7840 13132 7892 13184
rect 11060 13132 11112 13184
rect 11520 13132 11572 13184
rect 13084 13132 13136 13184
rect 20996 13268 21048 13320
rect 23756 13268 23808 13320
rect 24124 13311 24176 13320
rect 24124 13277 24133 13311
rect 24133 13277 24167 13311
rect 24167 13277 24176 13311
rect 24124 13268 24176 13277
rect 31852 13311 31904 13320
rect 31852 13277 31861 13311
rect 31861 13277 31895 13311
rect 31895 13277 31904 13311
rect 31852 13268 31904 13277
rect 32128 13311 32180 13320
rect 32128 13277 32137 13311
rect 32137 13277 32171 13311
rect 32171 13277 32180 13311
rect 32128 13268 32180 13277
rect 22468 13200 22520 13252
rect 33232 13200 33284 13252
rect 20904 13132 20956 13184
rect 21732 13132 21784 13184
rect 24032 13175 24084 13184
rect 24032 13141 24041 13175
rect 24041 13141 24075 13175
rect 24075 13141 24084 13175
rect 24032 13132 24084 13141
rect 28080 13132 28132 13184
rect 30472 13132 30524 13184
rect 6517 13030 6569 13082
rect 6581 13030 6633 13082
rect 6645 13030 6697 13082
rect 6709 13030 6761 13082
rect 17588 13030 17640 13082
rect 17652 13030 17704 13082
rect 17716 13030 17768 13082
rect 17780 13030 17832 13082
rect 28658 13030 28710 13082
rect 28722 13030 28774 13082
rect 28786 13030 28838 13082
rect 28850 13030 28902 13082
rect 2964 12928 3016 12980
rect 5448 12928 5500 12980
rect 8668 12971 8720 12980
rect 8668 12937 8677 12971
rect 8677 12937 8711 12971
rect 8711 12937 8720 12971
rect 8668 12928 8720 12937
rect 12624 12971 12676 12980
rect 12624 12937 12633 12971
rect 12633 12937 12667 12971
rect 12667 12937 12676 12971
rect 12624 12928 12676 12937
rect 14004 12971 14056 12980
rect 14004 12937 14013 12971
rect 14013 12937 14047 12971
rect 14047 12937 14056 12971
rect 14004 12928 14056 12937
rect 16304 12971 16356 12980
rect 16304 12937 16313 12971
rect 16313 12937 16347 12971
rect 16347 12937 16356 12971
rect 16304 12928 16356 12937
rect 20904 12928 20956 12980
rect 21272 12928 21324 12980
rect 21916 12928 21968 12980
rect 25044 12928 25096 12980
rect 26056 12971 26108 12980
rect 26056 12937 26065 12971
rect 26065 12937 26099 12971
rect 26099 12937 26108 12971
rect 26056 12928 26108 12937
rect 29552 12971 29604 12980
rect 29552 12937 29561 12971
rect 29561 12937 29595 12971
rect 29595 12937 29604 12971
rect 29552 12928 29604 12937
rect 30932 12928 30984 12980
rect 32128 12928 32180 12980
rect 1768 12835 1820 12844
rect 1768 12801 1777 12835
rect 1777 12801 1811 12835
rect 1811 12801 1820 12835
rect 1768 12792 1820 12801
rect 4712 12835 4764 12844
rect 4712 12801 4721 12835
rect 4721 12801 4755 12835
rect 4755 12801 4764 12835
rect 4712 12792 4764 12801
rect 7932 12835 7984 12844
rect 7932 12801 7941 12835
rect 7941 12801 7975 12835
rect 7975 12801 7984 12835
rect 7932 12792 7984 12801
rect 9588 12860 9640 12912
rect 10784 12860 10836 12912
rect 9128 12835 9180 12844
rect 9128 12801 9137 12835
rect 9137 12801 9171 12835
rect 9171 12801 9180 12835
rect 9128 12792 9180 12801
rect 11060 12792 11112 12844
rect 13636 12860 13688 12912
rect 12900 12792 12952 12844
rect 13176 12835 13228 12844
rect 13176 12801 13185 12835
rect 13185 12801 13219 12835
rect 13219 12801 13228 12835
rect 13176 12792 13228 12801
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 4068 12724 4120 12776
rect 7840 12767 7892 12776
rect 7840 12733 7849 12767
rect 7849 12733 7883 12767
rect 7883 12733 7892 12767
rect 7840 12724 7892 12733
rect 8760 12724 8812 12776
rect 12348 12724 12400 12776
rect 12808 12724 12860 12776
rect 13912 12724 13964 12776
rect 18788 12860 18840 12912
rect 19984 12860 20036 12912
rect 20720 12860 20772 12912
rect 22008 12860 22060 12912
rect 22468 12860 22520 12912
rect 26148 12903 26200 12912
rect 26148 12869 26157 12903
rect 26157 12869 26191 12903
rect 26191 12869 26200 12903
rect 26148 12860 26200 12869
rect 17960 12792 18012 12844
rect 23572 12792 23624 12844
rect 24032 12835 24084 12844
rect 24032 12801 24041 12835
rect 24041 12801 24075 12835
rect 24075 12801 24084 12835
rect 24032 12792 24084 12801
rect 26240 12835 26292 12844
rect 26240 12801 26249 12835
rect 26249 12801 26283 12835
rect 26283 12801 26292 12835
rect 26240 12792 26292 12801
rect 27620 12792 27672 12844
rect 27804 12835 27856 12844
rect 27804 12801 27813 12835
rect 27813 12801 27847 12835
rect 27847 12801 27856 12835
rect 27804 12792 27856 12801
rect 28080 12835 28132 12844
rect 28080 12801 28089 12835
rect 28089 12801 28123 12835
rect 28123 12801 28132 12835
rect 28080 12792 28132 12801
rect 30380 12903 30432 12912
rect 30380 12869 30389 12903
rect 30389 12869 30423 12903
rect 30423 12869 30432 12903
rect 30380 12860 30432 12869
rect 16212 12767 16264 12776
rect 16212 12733 16221 12767
rect 16221 12733 16255 12767
rect 16255 12733 16264 12767
rect 16212 12724 16264 12733
rect 17684 12767 17736 12776
rect 2688 12588 2740 12640
rect 5356 12656 5408 12708
rect 6000 12656 6052 12708
rect 5448 12588 5500 12640
rect 7104 12588 7156 12640
rect 14648 12588 14700 12640
rect 17684 12733 17693 12767
rect 17693 12733 17727 12767
rect 17727 12733 17736 12767
rect 17684 12724 17736 12733
rect 18052 12767 18104 12776
rect 18052 12733 18061 12767
rect 18061 12733 18095 12767
rect 18095 12733 18104 12767
rect 18052 12724 18104 12733
rect 18512 12767 18564 12776
rect 18512 12733 18521 12767
rect 18521 12733 18555 12767
rect 18555 12733 18564 12767
rect 18512 12724 18564 12733
rect 17960 12656 18012 12708
rect 22652 12724 22704 12776
rect 22376 12656 22428 12708
rect 23020 12724 23072 12776
rect 25964 12767 26016 12776
rect 25964 12733 25973 12767
rect 25973 12733 26007 12767
rect 26007 12733 26016 12767
rect 25964 12724 26016 12733
rect 29552 12724 29604 12776
rect 25044 12656 25096 12708
rect 28540 12656 28592 12708
rect 30472 12767 30524 12776
rect 30472 12733 30481 12767
rect 30481 12733 30515 12767
rect 30515 12733 30524 12767
rect 30472 12724 30524 12733
rect 31116 12767 31168 12776
rect 31116 12733 31125 12767
rect 31125 12733 31159 12767
rect 31159 12733 31168 12767
rect 31116 12724 31168 12733
rect 31760 12724 31812 12776
rect 33324 12767 33376 12776
rect 33324 12733 33333 12767
rect 33333 12733 33367 12767
rect 33367 12733 33376 12767
rect 33324 12724 33376 12733
rect 30288 12656 30340 12708
rect 30656 12656 30708 12708
rect 31300 12699 31352 12708
rect 31300 12665 31309 12699
rect 31309 12665 31343 12699
rect 31343 12665 31352 12699
rect 31300 12656 31352 12665
rect 33416 12656 33468 12708
rect 22744 12588 22796 12640
rect 24860 12588 24912 12640
rect 12052 12486 12104 12538
rect 12116 12486 12168 12538
rect 12180 12486 12232 12538
rect 12244 12486 12296 12538
rect 23123 12486 23175 12538
rect 23187 12486 23239 12538
rect 23251 12486 23303 12538
rect 23315 12486 23367 12538
rect 2872 12384 2924 12436
rect 7932 12384 7984 12436
rect 17684 12427 17736 12436
rect 17684 12393 17693 12427
rect 17693 12393 17727 12427
rect 17727 12393 17736 12427
rect 17684 12384 17736 12393
rect 17960 12384 18012 12436
rect 18236 12384 18288 12436
rect 21916 12384 21968 12436
rect 23020 12384 23072 12436
rect 23572 12427 23624 12436
rect 23572 12393 23581 12427
rect 23581 12393 23615 12427
rect 23615 12393 23624 12427
rect 23572 12384 23624 12393
rect 24124 12427 24176 12436
rect 24124 12393 24133 12427
rect 24133 12393 24167 12427
rect 24167 12393 24176 12427
rect 24124 12384 24176 12393
rect 1768 12359 1820 12368
rect 1768 12325 1777 12359
rect 1777 12325 1811 12359
rect 1811 12325 1820 12359
rect 1768 12316 1820 12325
rect 3884 12316 3936 12368
rect 5356 12316 5408 12368
rect 18144 12316 18196 12368
rect 4068 12248 4120 12300
rect 2964 12180 3016 12232
rect 3240 12180 3292 12232
rect 3976 12180 4028 12232
rect 4988 12223 5040 12232
rect 4988 12189 4997 12223
rect 4997 12189 5031 12223
rect 5031 12189 5040 12223
rect 4988 12180 5040 12189
rect 9864 12291 9916 12300
rect 9864 12257 9873 12291
rect 9873 12257 9907 12291
rect 9907 12257 9916 12291
rect 9864 12248 9916 12257
rect 13084 12291 13136 12300
rect 13084 12257 13093 12291
rect 13093 12257 13127 12291
rect 13127 12257 13136 12291
rect 13084 12248 13136 12257
rect 13452 12248 13504 12300
rect 16764 12291 16816 12300
rect 16764 12257 16773 12291
rect 16773 12257 16807 12291
rect 16807 12257 16816 12291
rect 16764 12248 16816 12257
rect 6000 12180 6052 12232
rect 9956 12223 10008 12232
rect 9956 12189 9965 12223
rect 9965 12189 9999 12223
rect 9999 12189 10008 12223
rect 9956 12180 10008 12189
rect 10048 12223 10100 12232
rect 10048 12189 10057 12223
rect 10057 12189 10091 12223
rect 10091 12189 10100 12223
rect 10048 12180 10100 12189
rect 15752 12180 15804 12232
rect 17316 12248 17368 12300
rect 17960 12248 18012 12300
rect 18880 12316 18932 12368
rect 20076 12316 20128 12368
rect 22008 12316 22060 12368
rect 22744 12359 22796 12368
rect 22744 12325 22753 12359
rect 22753 12325 22787 12359
rect 22787 12325 22796 12359
rect 22744 12316 22796 12325
rect 20168 12291 20220 12300
rect 20168 12257 20177 12291
rect 20177 12257 20211 12291
rect 20211 12257 20220 12291
rect 20168 12248 20220 12257
rect 23112 12316 23164 12368
rect 22652 12180 22704 12232
rect 23112 12180 23164 12232
rect 17224 12112 17276 12164
rect 20444 12112 20496 12164
rect 5448 12044 5500 12096
rect 8484 12087 8536 12096
rect 8484 12053 8493 12087
rect 8493 12053 8527 12087
rect 8527 12053 8536 12087
rect 8484 12044 8536 12053
rect 13268 12087 13320 12096
rect 13268 12053 13277 12087
rect 13277 12053 13311 12087
rect 13311 12053 13320 12087
rect 13268 12044 13320 12053
rect 15476 12087 15528 12096
rect 15476 12053 15485 12087
rect 15485 12053 15519 12087
rect 15519 12053 15528 12087
rect 15476 12044 15528 12053
rect 15568 12087 15620 12096
rect 15568 12053 15577 12087
rect 15577 12053 15611 12087
rect 15611 12053 15620 12087
rect 15568 12044 15620 12053
rect 18328 12044 18380 12096
rect 18788 12044 18840 12096
rect 19064 12044 19116 12096
rect 21364 12044 21416 12096
rect 25964 12384 26016 12436
rect 26148 12316 26200 12368
rect 28264 12384 28316 12436
rect 28540 12384 28592 12436
rect 29552 12427 29604 12436
rect 29552 12393 29561 12427
rect 29561 12393 29595 12427
rect 29595 12393 29604 12427
rect 29552 12384 29604 12393
rect 32496 12384 32548 12436
rect 24860 12248 24912 12300
rect 25596 12223 25648 12232
rect 25596 12189 25605 12223
rect 25605 12189 25639 12223
rect 25639 12189 25648 12223
rect 25596 12180 25648 12189
rect 25872 12180 25924 12232
rect 30380 12316 30432 12368
rect 33140 12316 33192 12368
rect 29460 12248 29512 12300
rect 30288 12248 30340 12300
rect 30748 12291 30800 12300
rect 30748 12257 30757 12291
rect 30757 12257 30791 12291
rect 30791 12257 30800 12291
rect 30748 12248 30800 12257
rect 31024 12291 31076 12300
rect 31024 12257 31033 12291
rect 31033 12257 31067 12291
rect 31067 12257 31076 12291
rect 31024 12248 31076 12257
rect 31116 12291 31168 12300
rect 31116 12257 31125 12291
rect 31125 12257 31159 12291
rect 31159 12257 31168 12291
rect 31116 12248 31168 12257
rect 31944 12248 31996 12300
rect 33508 12384 33560 12436
rect 33600 12359 33652 12368
rect 33600 12325 33609 12359
rect 33609 12325 33643 12359
rect 33643 12325 33652 12359
rect 33600 12316 33652 12325
rect 32956 12180 33008 12232
rect 26884 12112 26936 12164
rect 26608 12044 26660 12096
rect 32128 12087 32180 12096
rect 32128 12053 32137 12087
rect 32137 12053 32171 12087
rect 32171 12053 32180 12087
rect 32128 12044 32180 12053
rect 6517 11942 6569 11994
rect 6581 11942 6633 11994
rect 6645 11942 6697 11994
rect 6709 11942 6761 11994
rect 17588 11942 17640 11994
rect 17652 11942 17704 11994
rect 17716 11942 17768 11994
rect 17780 11942 17832 11994
rect 28658 11942 28710 11994
rect 28722 11942 28774 11994
rect 28786 11942 28838 11994
rect 28850 11942 28902 11994
rect 4988 11883 5040 11892
rect 4988 11849 4997 11883
rect 4997 11849 5031 11883
rect 5031 11849 5040 11883
rect 4988 11840 5040 11849
rect 9128 11883 9180 11892
rect 9128 11849 9137 11883
rect 9137 11849 9171 11883
rect 9171 11849 9180 11883
rect 9128 11840 9180 11849
rect 9864 11840 9916 11892
rect 12808 11840 12860 11892
rect 15200 11840 15252 11892
rect 2964 11772 3016 11824
rect 9956 11772 10008 11824
rect 10048 11772 10100 11824
rect 5448 11747 5500 11756
rect 5448 11713 5457 11747
rect 5457 11713 5491 11747
rect 5491 11713 5500 11747
rect 5448 11704 5500 11713
rect 3056 11636 3108 11688
rect 3424 11679 3476 11688
rect 3424 11645 3433 11679
rect 3433 11645 3467 11679
rect 3467 11645 3476 11679
rect 3424 11636 3476 11645
rect 5172 11636 5224 11688
rect 6000 11704 6052 11756
rect 7104 11747 7156 11756
rect 7104 11713 7113 11747
rect 7113 11713 7147 11747
rect 7147 11713 7156 11747
rect 7104 11704 7156 11713
rect 8484 11636 8536 11688
rect 10048 11636 10100 11688
rect 13636 11704 13688 11756
rect 16764 11840 16816 11892
rect 19248 11840 19300 11892
rect 20168 11840 20220 11892
rect 20444 11840 20496 11892
rect 25872 11840 25924 11892
rect 26240 11840 26292 11892
rect 32312 11772 32364 11824
rect 33232 11772 33284 11824
rect 16120 11704 16172 11756
rect 25596 11704 25648 11756
rect 27896 11704 27948 11756
rect 31392 11747 31444 11756
rect 31392 11713 31401 11747
rect 31401 11713 31435 11747
rect 31435 11713 31444 11747
rect 31392 11704 31444 11713
rect 10692 11636 10744 11688
rect 5540 11568 5592 11620
rect 9772 11568 9824 11620
rect 1768 11500 1820 11552
rect 8024 11500 8076 11552
rect 9680 11500 9732 11552
rect 10876 11500 10928 11552
rect 15568 11679 15620 11688
rect 15568 11645 15586 11679
rect 15586 11645 15620 11679
rect 15568 11636 15620 11645
rect 18512 11636 18564 11688
rect 14372 11568 14424 11620
rect 19064 11636 19116 11688
rect 24860 11636 24912 11688
rect 25044 11679 25096 11688
rect 25044 11645 25053 11679
rect 25053 11645 25087 11679
rect 25087 11645 25096 11679
rect 25044 11636 25096 11645
rect 25964 11636 26016 11688
rect 26608 11679 26660 11688
rect 26608 11645 26617 11679
rect 26617 11645 26651 11679
rect 26651 11645 26660 11679
rect 26608 11636 26660 11645
rect 28172 11679 28224 11688
rect 28172 11645 28181 11679
rect 28181 11645 28215 11679
rect 28215 11645 28224 11679
rect 28172 11636 28224 11645
rect 28448 11679 28500 11688
rect 28448 11645 28457 11679
rect 28457 11645 28491 11679
rect 28491 11645 28500 11679
rect 28448 11636 28500 11645
rect 29552 11679 29604 11688
rect 29552 11645 29561 11679
rect 29561 11645 29595 11679
rect 29595 11645 29604 11679
rect 29552 11636 29604 11645
rect 30380 11636 30432 11688
rect 30748 11679 30800 11688
rect 30748 11645 30757 11679
rect 30757 11645 30791 11679
rect 30791 11645 30800 11679
rect 30748 11636 30800 11645
rect 31024 11636 31076 11688
rect 31300 11636 31352 11688
rect 33232 11636 33284 11688
rect 21272 11568 21324 11620
rect 28264 11568 28316 11620
rect 11796 11500 11848 11552
rect 13084 11500 13136 11552
rect 13728 11500 13780 11552
rect 14464 11543 14516 11552
rect 14464 11509 14473 11543
rect 14473 11509 14507 11543
rect 14507 11509 14516 11543
rect 14464 11500 14516 11509
rect 23572 11500 23624 11552
rect 27804 11500 27856 11552
rect 33324 11543 33376 11552
rect 33324 11509 33333 11543
rect 33333 11509 33367 11543
rect 33367 11509 33376 11543
rect 33324 11500 33376 11509
rect 12052 11398 12104 11450
rect 12116 11398 12168 11450
rect 12180 11398 12232 11450
rect 12244 11398 12296 11450
rect 23123 11398 23175 11450
rect 23187 11398 23239 11450
rect 23251 11398 23303 11450
rect 23315 11398 23367 11450
rect 9772 11296 9824 11348
rect 2688 11228 2740 11280
rect 9680 11271 9732 11280
rect 9680 11237 9689 11271
rect 9689 11237 9723 11271
rect 9723 11237 9732 11271
rect 9680 11228 9732 11237
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 1768 11203 1820 11212
rect 1768 11169 1777 11203
rect 1777 11169 1811 11203
rect 1811 11169 1820 11203
rect 1768 11160 1820 11169
rect 5264 11203 5316 11212
rect 5264 11169 5273 11203
rect 5273 11169 5307 11203
rect 5307 11169 5316 11203
rect 5264 11160 5316 11169
rect 5540 11160 5592 11212
rect 10784 11228 10836 11280
rect 11152 11228 11204 11280
rect 13268 11296 13320 11348
rect 15752 11339 15804 11348
rect 15752 11305 15761 11339
rect 15761 11305 15795 11339
rect 15795 11305 15804 11339
rect 15752 11296 15804 11305
rect 18052 11339 18104 11348
rect 18052 11305 18061 11339
rect 18061 11305 18095 11339
rect 18095 11305 18104 11339
rect 18052 11296 18104 11305
rect 19984 11296 20036 11348
rect 23020 11296 23072 11348
rect 31024 11296 31076 11348
rect 2872 11092 2924 11144
rect 3056 11092 3108 11144
rect 5172 11092 5224 11144
rect 10692 11092 10744 11144
rect 13452 11160 13504 11212
rect 13728 11203 13780 11212
rect 13728 11169 13737 11203
rect 13737 11169 13771 11203
rect 13771 11169 13780 11203
rect 13728 11160 13780 11169
rect 13268 11024 13320 11076
rect 14096 11228 14148 11280
rect 14464 11160 14516 11212
rect 15844 11203 15896 11212
rect 15844 11169 15853 11203
rect 15853 11169 15887 11203
rect 15887 11169 15896 11203
rect 15844 11160 15896 11169
rect 18512 11228 18564 11280
rect 26884 11228 26936 11280
rect 27804 11271 27856 11280
rect 27804 11237 27813 11271
rect 27813 11237 27847 11271
rect 27847 11237 27856 11271
rect 27804 11228 27856 11237
rect 28264 11228 28316 11280
rect 32128 11271 32180 11280
rect 32128 11237 32137 11271
rect 32137 11237 32171 11271
rect 32171 11237 32180 11271
rect 32128 11228 32180 11237
rect 32588 11228 32640 11280
rect 18144 11160 18196 11212
rect 19800 11160 19852 11212
rect 20352 11160 20404 11212
rect 21732 11203 21784 11212
rect 21732 11169 21741 11203
rect 21741 11169 21775 11203
rect 21775 11169 21784 11203
rect 21732 11160 21784 11169
rect 22376 11203 22428 11212
rect 22376 11169 22385 11203
rect 22385 11169 22419 11203
rect 22419 11169 22428 11203
rect 22376 11160 22428 11169
rect 22560 11203 22612 11212
rect 22560 11169 22569 11203
rect 22569 11169 22603 11203
rect 22603 11169 22612 11203
rect 22560 11160 22612 11169
rect 22836 11160 22888 11212
rect 23572 11203 23624 11212
rect 23572 11169 23581 11203
rect 23581 11169 23615 11203
rect 23615 11169 23624 11203
rect 23572 11160 23624 11169
rect 25688 11160 25740 11212
rect 19248 11092 19300 11144
rect 23848 11135 23900 11144
rect 23848 11101 23857 11135
rect 23857 11101 23891 11135
rect 23891 11101 23900 11135
rect 23848 11092 23900 11101
rect 25964 11092 26016 11144
rect 26608 11160 26660 11212
rect 27896 11092 27948 11144
rect 29092 11092 29144 11144
rect 31208 11160 31260 11212
rect 31852 11203 31904 11212
rect 31852 11169 31861 11203
rect 31861 11169 31895 11203
rect 31895 11169 31904 11203
rect 31852 11160 31904 11169
rect 14188 11024 14240 11076
rect 18420 11024 18472 11076
rect 18972 11067 19024 11076
rect 18972 11033 18981 11067
rect 18981 11033 19015 11067
rect 19015 11033 19024 11067
rect 18972 11024 19024 11033
rect 21548 11024 21600 11076
rect 21916 11024 21968 11076
rect 23480 11024 23532 11076
rect 26976 11067 27028 11076
rect 26976 11033 26985 11067
rect 26985 11033 27019 11067
rect 27019 11033 27028 11067
rect 26976 11024 27028 11033
rect 2780 10956 2832 11008
rect 3424 10956 3476 11008
rect 4896 10999 4948 11008
rect 4896 10965 4905 10999
rect 4905 10965 4939 10999
rect 4939 10965 4948 10999
rect 4896 10956 4948 10965
rect 10416 10956 10468 11008
rect 14924 10999 14976 11008
rect 14924 10965 14933 10999
rect 14933 10965 14967 10999
rect 14967 10965 14976 10999
rect 14924 10956 14976 10965
rect 17224 10999 17276 11008
rect 17224 10965 17233 10999
rect 17233 10965 17267 10999
rect 17267 10965 17276 10999
rect 17224 10956 17276 10965
rect 17408 10999 17460 11008
rect 17408 10965 17417 10999
rect 17417 10965 17451 10999
rect 17451 10965 17460 10999
rect 17408 10956 17460 10965
rect 23756 10999 23808 11008
rect 23756 10965 23765 10999
rect 23765 10965 23799 10999
rect 23799 10965 23808 10999
rect 23756 10956 23808 10965
rect 25412 10956 25464 11008
rect 28448 10956 28500 11008
rect 29644 10956 29696 11008
rect 30656 10956 30708 11008
rect 33232 10956 33284 11008
rect 6517 10854 6569 10906
rect 6581 10854 6633 10906
rect 6645 10854 6697 10906
rect 6709 10854 6761 10906
rect 17588 10854 17640 10906
rect 17652 10854 17704 10906
rect 17716 10854 17768 10906
rect 17780 10854 17832 10906
rect 28658 10854 28710 10906
rect 28722 10854 28774 10906
rect 28786 10854 28838 10906
rect 28850 10854 28902 10906
rect 3056 10752 3108 10804
rect 5540 10752 5592 10804
rect 10048 10752 10100 10804
rect 10416 10795 10468 10804
rect 10416 10761 10425 10795
rect 10425 10761 10459 10795
rect 10459 10761 10468 10795
rect 10416 10752 10468 10761
rect 12348 10752 12400 10804
rect 13360 10795 13412 10804
rect 13360 10761 13369 10795
rect 13369 10761 13403 10795
rect 13403 10761 13412 10795
rect 13360 10752 13412 10761
rect 14372 10795 14424 10804
rect 14372 10761 14381 10795
rect 14381 10761 14415 10795
rect 14415 10761 14424 10795
rect 14372 10752 14424 10761
rect 15476 10752 15528 10804
rect 16396 10752 16448 10804
rect 18328 10752 18380 10804
rect 19800 10795 19852 10804
rect 19800 10761 19809 10795
rect 19809 10761 19843 10795
rect 19843 10761 19852 10795
rect 19800 10752 19852 10761
rect 16488 10684 16540 10736
rect 2872 10616 2924 10668
rect 3976 10659 4028 10668
rect 3976 10625 3985 10659
rect 3985 10625 4019 10659
rect 4019 10625 4028 10659
rect 3976 10616 4028 10625
rect 4896 10616 4948 10668
rect 8852 10659 8904 10668
rect 8852 10625 8861 10659
rect 8861 10625 8895 10659
rect 8895 10625 8904 10659
rect 8852 10616 8904 10625
rect 9588 10616 9640 10668
rect 3332 10548 3384 10600
rect 8300 10548 8352 10600
rect 9864 10548 9916 10600
rect 10876 10548 10928 10600
rect 11060 10548 11112 10600
rect 11520 10548 11572 10600
rect 11888 10548 11940 10600
rect 13544 10616 13596 10668
rect 14924 10616 14976 10668
rect 15660 10616 15712 10668
rect 13268 10591 13320 10600
rect 13268 10557 13277 10591
rect 13277 10557 13311 10591
rect 13311 10557 13320 10591
rect 13268 10548 13320 10557
rect 5356 10480 5408 10532
rect 8576 10523 8628 10532
rect 8576 10489 8585 10523
rect 8585 10489 8619 10523
rect 8619 10489 8628 10523
rect 8576 10480 8628 10489
rect 13176 10480 13228 10532
rect 13728 10548 13780 10600
rect 14188 10591 14240 10600
rect 14188 10557 14197 10591
rect 14197 10557 14231 10591
rect 14231 10557 14240 10591
rect 14188 10548 14240 10557
rect 15200 10591 15252 10600
rect 15200 10557 15209 10591
rect 15209 10557 15243 10591
rect 15243 10557 15252 10591
rect 15200 10548 15252 10557
rect 18420 10616 18472 10668
rect 18604 10659 18656 10668
rect 18604 10625 18613 10659
rect 18613 10625 18647 10659
rect 18647 10625 18656 10659
rect 18604 10616 18656 10625
rect 14096 10480 14148 10532
rect 8208 10455 8260 10464
rect 8208 10421 8217 10455
rect 8217 10421 8251 10455
rect 8251 10421 8260 10455
rect 8208 10412 8260 10421
rect 8668 10455 8720 10464
rect 8668 10421 8677 10455
rect 8677 10421 8711 10455
rect 8711 10421 8720 10455
rect 8668 10412 8720 10421
rect 10232 10412 10284 10464
rect 11060 10412 11112 10464
rect 13268 10412 13320 10464
rect 15476 10455 15528 10464
rect 15476 10421 15485 10455
rect 15485 10421 15519 10455
rect 15519 10421 15528 10455
rect 15476 10412 15528 10421
rect 17224 10548 17276 10600
rect 18236 10591 18288 10600
rect 18236 10557 18245 10591
rect 18245 10557 18279 10591
rect 18279 10557 18288 10591
rect 18236 10548 18288 10557
rect 19248 10591 19300 10600
rect 18144 10480 18196 10532
rect 19248 10557 19257 10591
rect 19257 10557 19291 10591
rect 19291 10557 19300 10591
rect 19248 10548 19300 10557
rect 19984 10480 20036 10532
rect 16396 10412 16448 10464
rect 20812 10412 20864 10464
rect 21272 10616 21324 10668
rect 24584 10616 24636 10668
rect 25596 10752 25648 10804
rect 26884 10795 26936 10804
rect 26884 10761 26893 10795
rect 26893 10761 26927 10795
rect 26927 10761 26936 10795
rect 26884 10752 26936 10761
rect 29552 10752 29604 10804
rect 29644 10752 29696 10804
rect 33140 10795 33192 10804
rect 33140 10761 33149 10795
rect 33149 10761 33183 10795
rect 33183 10761 33192 10795
rect 33140 10752 33192 10761
rect 31208 10684 31260 10736
rect 25412 10659 25464 10668
rect 25412 10625 25421 10659
rect 25421 10625 25455 10659
rect 25455 10625 25464 10659
rect 25412 10616 25464 10625
rect 29644 10616 29696 10668
rect 30380 10616 30432 10668
rect 23756 10548 23808 10600
rect 29092 10591 29144 10600
rect 29092 10557 29101 10591
rect 29101 10557 29135 10591
rect 29135 10557 29144 10591
rect 29092 10548 29144 10557
rect 30656 10591 30708 10600
rect 27160 10480 27212 10532
rect 28264 10480 28316 10532
rect 23020 10455 23072 10464
rect 23020 10421 23029 10455
rect 23029 10421 23063 10455
rect 23063 10421 23072 10455
rect 23020 10412 23072 10421
rect 30656 10557 30665 10591
rect 30665 10557 30699 10591
rect 30699 10557 30708 10591
rect 30656 10548 30708 10557
rect 31024 10616 31076 10668
rect 31484 10548 31536 10600
rect 33416 10616 33468 10668
rect 33232 10591 33284 10600
rect 33232 10557 33241 10591
rect 33241 10557 33275 10591
rect 33275 10557 33284 10591
rect 33232 10548 33284 10557
rect 31668 10480 31720 10532
rect 31300 10412 31352 10464
rect 12052 10310 12104 10362
rect 12116 10310 12168 10362
rect 12180 10310 12232 10362
rect 12244 10310 12296 10362
rect 23123 10310 23175 10362
rect 23187 10310 23239 10362
rect 23251 10310 23303 10362
rect 23315 10310 23367 10362
rect 2780 10251 2832 10260
rect 2780 10217 2789 10251
rect 2789 10217 2823 10251
rect 2823 10217 2832 10251
rect 10232 10251 10284 10260
rect 2780 10208 2832 10217
rect 10232 10217 10241 10251
rect 10241 10217 10275 10251
rect 10275 10217 10284 10251
rect 10232 10208 10284 10217
rect 13268 10251 13320 10260
rect 13268 10217 13277 10251
rect 13277 10217 13311 10251
rect 13311 10217 13320 10251
rect 13268 10208 13320 10217
rect 14740 10251 14792 10260
rect 14740 10217 14749 10251
rect 14749 10217 14783 10251
rect 14783 10217 14792 10251
rect 14740 10208 14792 10217
rect 15568 10208 15620 10260
rect 16488 10208 16540 10260
rect 19984 10251 20036 10260
rect 9312 10140 9364 10192
rect 8208 10115 8260 10124
rect 8208 10081 8217 10115
rect 8217 10081 8251 10115
rect 8251 10081 8260 10115
rect 8208 10072 8260 10081
rect 8760 10072 8812 10124
rect 9404 10072 9456 10124
rect 12808 10140 12860 10192
rect 15476 10140 15528 10192
rect 16764 10140 16816 10192
rect 17316 10140 17368 10192
rect 11336 10115 11388 10124
rect 2872 10047 2924 10056
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 3332 10004 3384 10056
rect 8116 10004 8168 10056
rect 10140 10004 10192 10056
rect 8392 9936 8444 9988
rect 11336 10081 11345 10115
rect 11345 10081 11379 10115
rect 11379 10081 11388 10115
rect 11336 10072 11388 10081
rect 13452 10115 13504 10124
rect 11428 10047 11480 10056
rect 11428 10013 11437 10047
rect 11437 10013 11471 10047
rect 11471 10013 11480 10047
rect 11428 10004 11480 10013
rect 11520 10047 11572 10056
rect 11520 10013 11529 10047
rect 11529 10013 11563 10047
rect 11563 10013 11572 10047
rect 11520 10004 11572 10013
rect 1768 9868 1820 9920
rect 7104 9868 7156 9920
rect 9680 9868 9732 9920
rect 11888 9868 11940 9920
rect 13452 10081 13461 10115
rect 13461 10081 13495 10115
rect 13495 10081 13504 10115
rect 13452 10072 13504 10081
rect 16120 10115 16172 10124
rect 16120 10081 16129 10115
rect 16129 10081 16163 10115
rect 16163 10081 16172 10115
rect 16120 10072 16172 10081
rect 16672 10115 16724 10124
rect 16672 10081 16681 10115
rect 16681 10081 16715 10115
rect 16715 10081 16724 10115
rect 16672 10072 16724 10081
rect 16948 10115 17000 10124
rect 16948 10081 16957 10115
rect 16957 10081 16991 10115
rect 16991 10081 17000 10115
rect 16948 10072 17000 10081
rect 17408 10115 17460 10124
rect 17408 10081 17417 10115
rect 17417 10081 17451 10115
rect 17451 10081 17460 10115
rect 17408 10072 17460 10081
rect 17960 10072 18012 10124
rect 19984 10217 19993 10251
rect 19993 10217 20027 10251
rect 20027 10217 20036 10251
rect 19984 10208 20036 10217
rect 22560 10208 22612 10260
rect 23848 10208 23900 10260
rect 29644 10208 29696 10260
rect 27160 10140 27212 10192
rect 30196 10140 30248 10192
rect 20812 10115 20864 10124
rect 17316 10004 17368 10056
rect 19984 10047 20036 10056
rect 19984 10013 19993 10047
rect 19993 10013 20027 10047
rect 20027 10013 20036 10047
rect 19984 10004 20036 10013
rect 20812 10081 20821 10115
rect 20821 10081 20855 10115
rect 20855 10081 20864 10115
rect 20812 10072 20864 10081
rect 21364 10072 21416 10124
rect 20536 10004 20588 10056
rect 17132 9868 17184 9920
rect 23020 10072 23072 10124
rect 22376 10004 22428 10056
rect 25596 10072 25648 10124
rect 30748 10115 30800 10124
rect 30748 10081 30757 10115
rect 30757 10081 30791 10115
rect 30791 10081 30800 10115
rect 30748 10072 30800 10081
rect 31116 10115 31168 10124
rect 29092 9936 29144 9988
rect 31116 10081 31125 10115
rect 31125 10081 31159 10115
rect 31159 10081 31168 10115
rect 31116 10072 31168 10081
rect 31484 10072 31536 10124
rect 32312 10140 32364 10192
rect 32404 10115 32456 10124
rect 31300 10004 31352 10056
rect 32404 10081 32413 10115
rect 32413 10081 32447 10115
rect 32447 10081 32456 10115
rect 32404 10072 32456 10081
rect 31668 9936 31720 9988
rect 33416 9936 33468 9988
rect 22836 9911 22888 9920
rect 22836 9877 22845 9911
rect 22845 9877 22879 9911
rect 22879 9877 22888 9911
rect 22836 9868 22888 9877
rect 28356 9911 28408 9920
rect 28356 9877 28365 9911
rect 28365 9877 28399 9911
rect 28399 9877 28408 9911
rect 28356 9868 28408 9877
rect 33140 9868 33192 9920
rect 33324 9911 33376 9920
rect 33324 9877 33333 9911
rect 33333 9877 33367 9911
rect 33367 9877 33376 9911
rect 33324 9868 33376 9877
rect 6517 9766 6569 9818
rect 6581 9766 6633 9818
rect 6645 9766 6697 9818
rect 6709 9766 6761 9818
rect 17588 9766 17640 9818
rect 17652 9766 17704 9818
rect 17716 9766 17768 9818
rect 17780 9766 17832 9818
rect 28658 9766 28710 9818
rect 28722 9766 28774 9818
rect 28786 9766 28838 9818
rect 28850 9766 28902 9818
rect 2872 9664 2924 9716
rect 8576 9664 8628 9716
rect 11336 9664 11388 9716
rect 15660 9707 15712 9716
rect 15660 9673 15669 9707
rect 15669 9673 15703 9707
rect 15703 9673 15712 9707
rect 15660 9664 15712 9673
rect 19984 9664 20036 9716
rect 21364 9707 21416 9716
rect 21364 9673 21373 9707
rect 21373 9673 21407 9707
rect 21407 9673 21416 9707
rect 21364 9664 21416 9673
rect 11060 9639 11112 9648
rect 11060 9605 11069 9639
rect 11069 9605 11103 9639
rect 11103 9605 11112 9639
rect 11060 9596 11112 9605
rect 16856 9596 16908 9648
rect 21180 9596 21232 9648
rect 25964 9639 26016 9648
rect 25964 9605 25973 9639
rect 25973 9605 26007 9639
rect 26007 9605 26016 9639
rect 25964 9596 26016 9605
rect 1768 9571 1820 9580
rect 1768 9537 1777 9571
rect 1777 9537 1811 9571
rect 1811 9537 1820 9571
rect 1768 9528 1820 9537
rect 5264 9528 5316 9580
rect 7104 9571 7156 9580
rect 1492 9460 1544 9512
rect 3792 9460 3844 9512
rect 4436 9460 4488 9512
rect 7104 9537 7113 9571
rect 7113 9537 7147 9571
rect 7147 9537 7156 9571
rect 7104 9528 7156 9537
rect 9220 9528 9272 9580
rect 9404 9528 9456 9580
rect 9772 9571 9824 9580
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 9772 9528 9824 9537
rect 12900 9528 12952 9580
rect 13360 9528 13412 9580
rect 13636 9528 13688 9580
rect 21916 9528 21968 9580
rect 24584 9571 24636 9580
rect 24584 9537 24593 9571
rect 24593 9537 24627 9571
rect 24627 9537 24636 9571
rect 24584 9528 24636 9537
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 8668 9460 8720 9512
rect 9496 9503 9548 9512
rect 9496 9469 9505 9503
rect 9505 9469 9539 9503
rect 9539 9469 9548 9503
rect 9496 9460 9548 9469
rect 2320 9392 2372 9444
rect 3332 9392 3384 9444
rect 5632 9392 5684 9444
rect 8116 9392 8168 9444
rect 8392 9392 8444 9444
rect 13452 9460 13504 9512
rect 15568 9503 15620 9512
rect 15568 9469 15577 9503
rect 15577 9469 15611 9503
rect 15611 9469 15620 9503
rect 15568 9460 15620 9469
rect 11428 9392 11480 9444
rect 15844 9460 15896 9512
rect 17316 9503 17368 9512
rect 17316 9469 17325 9503
rect 17325 9469 17359 9503
rect 17359 9469 17368 9503
rect 17316 9460 17368 9469
rect 18604 9460 18656 9512
rect 19800 9460 19852 9512
rect 20352 9460 20404 9512
rect 21548 9503 21600 9512
rect 21548 9469 21557 9503
rect 21557 9469 21591 9503
rect 21591 9469 21600 9503
rect 21548 9460 21600 9469
rect 22560 9503 22612 9512
rect 22560 9469 22569 9503
rect 22569 9469 22603 9503
rect 22603 9469 22612 9503
rect 22560 9460 22612 9469
rect 24400 9460 24452 9512
rect 29000 9503 29052 9512
rect 29000 9469 29009 9503
rect 29009 9469 29043 9503
rect 29043 9469 29052 9503
rect 29000 9460 29052 9469
rect 29460 9503 29512 9512
rect 29460 9469 29469 9503
rect 29469 9469 29503 9503
rect 29503 9469 29512 9503
rect 29460 9460 29512 9469
rect 29736 9503 29788 9512
rect 29736 9469 29745 9503
rect 29745 9469 29779 9503
rect 29779 9469 29788 9503
rect 29736 9460 29788 9469
rect 4620 9324 4672 9376
rect 9588 9367 9640 9376
rect 9588 9333 9597 9367
rect 9597 9333 9631 9367
rect 9631 9333 9640 9367
rect 12532 9367 12584 9376
rect 9588 9324 9640 9333
rect 12532 9333 12541 9367
rect 12541 9333 12575 9367
rect 12575 9333 12584 9367
rect 12532 9324 12584 9333
rect 20076 9392 20128 9444
rect 23572 9392 23624 9444
rect 33416 9664 33468 9716
rect 30748 9639 30800 9648
rect 30748 9605 30757 9639
rect 30757 9605 30791 9639
rect 30791 9605 30800 9639
rect 30748 9596 30800 9605
rect 30748 9460 30800 9512
rect 32404 9528 32456 9580
rect 31208 9503 31260 9512
rect 31208 9469 31217 9503
rect 31217 9469 31251 9503
rect 31251 9469 31260 9503
rect 31208 9460 31260 9469
rect 31300 9460 31352 9512
rect 13636 9367 13688 9376
rect 13636 9333 13645 9367
rect 13645 9333 13679 9367
rect 13679 9333 13688 9367
rect 13636 9324 13688 9333
rect 20628 9324 20680 9376
rect 20812 9367 20864 9376
rect 20812 9333 20821 9367
rect 20821 9333 20855 9367
rect 20855 9333 20864 9367
rect 20812 9324 20864 9333
rect 20904 9324 20956 9376
rect 23848 9324 23900 9376
rect 12052 9222 12104 9274
rect 12116 9222 12168 9274
rect 12180 9222 12232 9274
rect 12244 9222 12296 9274
rect 23123 9222 23175 9274
rect 23187 9222 23239 9274
rect 23251 9222 23303 9274
rect 23315 9222 23367 9274
rect 5264 9120 5316 9172
rect 9588 9120 9640 9172
rect 12532 9120 12584 9172
rect 5356 9052 5408 9104
rect 2872 8984 2924 9036
rect 4620 9027 4672 9036
rect 4620 8993 4629 9027
rect 4629 8993 4663 9027
rect 4663 8993 4672 9027
rect 4620 8984 4672 8993
rect 8392 9027 8444 9036
rect 8392 8993 8401 9027
rect 8401 8993 8435 9027
rect 8435 8993 8444 9027
rect 8392 8984 8444 8993
rect 9864 9052 9916 9104
rect 9680 9027 9732 9036
rect 2964 8916 3016 8968
rect 4528 8916 4580 8968
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 10232 8984 10284 9036
rect 9036 8916 9088 8968
rect 11060 8984 11112 9036
rect 11612 8984 11664 9036
rect 13452 9120 13504 9172
rect 13636 9163 13688 9172
rect 13636 9129 13645 9163
rect 13645 9129 13679 9163
rect 13679 9129 13688 9163
rect 13636 9120 13688 9129
rect 15200 9120 15252 9172
rect 16672 9120 16724 9172
rect 17224 9163 17276 9172
rect 17224 9129 17233 9163
rect 17233 9129 17267 9163
rect 17267 9129 17276 9163
rect 17224 9120 17276 9129
rect 18236 9163 18288 9172
rect 18236 9129 18245 9163
rect 18245 9129 18279 9163
rect 18279 9129 18288 9163
rect 18236 9120 18288 9129
rect 20352 9120 20404 9172
rect 12808 9027 12860 9036
rect 12808 8993 12817 9027
rect 12817 8993 12851 9027
rect 12851 8993 12860 9027
rect 12808 8984 12860 8993
rect 13268 9027 13320 9036
rect 13268 8993 13277 9027
rect 13277 8993 13311 9027
rect 13311 8993 13320 9027
rect 13268 8984 13320 8993
rect 16120 8984 16172 9036
rect 16212 8984 16264 9036
rect 17224 8984 17276 9036
rect 17960 8984 18012 9036
rect 20904 9052 20956 9104
rect 22376 9120 22428 9172
rect 23572 9163 23624 9172
rect 23572 9129 23581 9163
rect 23581 9129 23615 9163
rect 23615 9129 23624 9163
rect 23572 9120 23624 9129
rect 29092 9120 29144 9172
rect 29460 9163 29512 9172
rect 29460 9129 29469 9163
rect 29469 9129 29503 9163
rect 29503 9129 29512 9163
rect 29460 9120 29512 9129
rect 30748 9095 30800 9104
rect 30748 9061 30757 9095
rect 30757 9061 30791 9095
rect 30791 9061 30800 9095
rect 30748 9052 30800 9061
rect 33232 9120 33284 9172
rect 9496 8848 9548 8900
rect 19708 8916 19760 8968
rect 20812 8984 20864 9036
rect 23848 9027 23900 9036
rect 22100 8916 22152 8968
rect 23848 8993 23857 9027
rect 23857 8993 23891 9027
rect 23891 8993 23900 9027
rect 23848 8984 23900 8993
rect 27068 8984 27120 9036
rect 28356 8984 28408 9036
rect 30932 9027 30984 9036
rect 30932 8993 30941 9027
rect 30941 8993 30975 9027
rect 30975 8993 30984 9027
rect 30932 8984 30984 8993
rect 32588 9052 32640 9104
rect 23572 8959 23624 8968
rect 23572 8925 23581 8959
rect 23581 8925 23615 8959
rect 23615 8925 23624 8959
rect 23572 8916 23624 8925
rect 25964 8959 26016 8968
rect 3148 8780 3200 8832
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 20168 8848 20220 8900
rect 20536 8891 20588 8900
rect 20536 8857 20545 8891
rect 20545 8857 20579 8891
rect 20579 8857 20588 8891
rect 20536 8848 20588 8857
rect 21180 8848 21232 8900
rect 23480 8848 23532 8900
rect 23848 8848 23900 8900
rect 18880 8823 18932 8832
rect 18880 8789 18889 8823
rect 18889 8789 18923 8823
rect 18923 8789 18932 8823
rect 18880 8780 18932 8789
rect 18972 8823 19024 8832
rect 18972 8789 18981 8823
rect 18981 8789 19015 8823
rect 19015 8789 19024 8823
rect 25964 8925 25973 8959
rect 25973 8925 26007 8959
rect 26007 8925 26016 8959
rect 25964 8916 26016 8925
rect 29092 8916 29144 8968
rect 31024 8916 31076 8968
rect 31852 8959 31904 8968
rect 31852 8925 31861 8959
rect 31861 8925 31895 8959
rect 31895 8925 31904 8959
rect 31852 8916 31904 8925
rect 32312 8916 32364 8968
rect 18972 8780 19024 8789
rect 26056 8780 26108 8832
rect 28172 8780 28224 8832
rect 28540 8823 28592 8832
rect 28540 8789 28549 8823
rect 28549 8789 28583 8823
rect 28583 8789 28592 8823
rect 28540 8780 28592 8789
rect 6517 8678 6569 8730
rect 6581 8678 6633 8730
rect 6645 8678 6697 8730
rect 6709 8678 6761 8730
rect 17588 8678 17640 8730
rect 17652 8678 17704 8730
rect 17716 8678 17768 8730
rect 17780 8678 17832 8730
rect 28658 8678 28710 8730
rect 28722 8678 28774 8730
rect 28786 8678 28838 8730
rect 28850 8678 28902 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 4436 8619 4488 8628
rect 4436 8585 4445 8619
rect 4445 8585 4479 8619
rect 4479 8585 4488 8619
rect 4436 8576 4488 8585
rect 5724 8576 5776 8628
rect 16212 8576 16264 8628
rect 16948 8576 17000 8628
rect 17132 8576 17184 8628
rect 17960 8576 18012 8628
rect 19800 8576 19852 8628
rect 20168 8576 20220 8628
rect 4528 8508 4580 8560
rect 6828 8508 6880 8560
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 3148 8415 3200 8424
rect 3148 8381 3157 8415
rect 3157 8381 3191 8415
rect 3191 8381 3200 8415
rect 3148 8372 3200 8381
rect 3792 8372 3844 8424
rect 8576 8347 8628 8356
rect 8576 8313 8585 8347
rect 8585 8313 8619 8347
rect 8619 8313 8628 8347
rect 8576 8304 8628 8313
rect 11336 8508 11388 8560
rect 25964 8576 26016 8628
rect 31852 8576 31904 8628
rect 9680 8440 9732 8492
rect 11520 8440 11572 8492
rect 20628 8440 20680 8492
rect 11888 8372 11940 8424
rect 15384 8415 15436 8424
rect 9772 8304 9824 8356
rect 10968 8304 11020 8356
rect 12900 8304 12952 8356
rect 15384 8381 15393 8415
rect 15393 8381 15427 8415
rect 15427 8381 15436 8415
rect 15384 8372 15436 8381
rect 16120 8372 16172 8424
rect 17040 8372 17092 8424
rect 17960 8415 18012 8424
rect 17960 8381 17969 8415
rect 17969 8381 18003 8415
rect 18003 8381 18012 8415
rect 17960 8372 18012 8381
rect 18696 8415 18748 8424
rect 18696 8381 18705 8415
rect 18705 8381 18739 8415
rect 18739 8381 18748 8415
rect 18696 8372 18748 8381
rect 18972 8415 19024 8424
rect 18972 8381 19006 8415
rect 19006 8381 19024 8415
rect 18972 8372 19024 8381
rect 22100 8372 22152 8424
rect 17224 8304 17276 8356
rect 18788 8304 18840 8356
rect 19156 8304 19208 8356
rect 22560 8347 22612 8356
rect 2780 8279 2832 8288
rect 2780 8245 2789 8279
rect 2789 8245 2823 8279
rect 2823 8245 2832 8279
rect 3240 8279 3292 8288
rect 2780 8236 2832 8245
rect 3240 8245 3249 8279
rect 3249 8245 3283 8279
rect 3283 8245 3292 8279
rect 3240 8236 3292 8245
rect 8208 8279 8260 8288
rect 8208 8245 8217 8279
rect 8217 8245 8251 8279
rect 8251 8245 8260 8279
rect 8208 8236 8260 8245
rect 8668 8279 8720 8288
rect 8668 8245 8677 8279
rect 8677 8245 8711 8279
rect 8711 8245 8720 8279
rect 8668 8236 8720 8245
rect 9956 8236 10008 8288
rect 10416 8279 10468 8288
rect 10416 8245 10425 8279
rect 10425 8245 10459 8279
rect 10459 8245 10468 8279
rect 10416 8236 10468 8245
rect 10784 8236 10836 8288
rect 12624 8279 12676 8288
rect 12624 8245 12633 8279
rect 12633 8245 12667 8279
rect 12667 8245 12676 8279
rect 12624 8236 12676 8245
rect 12992 8279 13044 8288
rect 12992 8245 13001 8279
rect 13001 8245 13035 8279
rect 13035 8245 13044 8279
rect 12992 8236 13044 8245
rect 13452 8236 13504 8288
rect 15568 8236 15620 8288
rect 22560 8313 22569 8347
rect 22569 8313 22603 8347
rect 22603 8313 22612 8347
rect 22560 8304 22612 8313
rect 22836 8372 22888 8424
rect 26056 8372 26108 8424
rect 28172 8415 28224 8424
rect 28172 8381 28181 8415
rect 28181 8381 28215 8415
rect 28215 8381 28224 8415
rect 28172 8372 28224 8381
rect 30472 8440 30524 8492
rect 30932 8440 30984 8492
rect 29920 8372 29972 8424
rect 30104 8415 30156 8424
rect 30104 8381 30113 8415
rect 30113 8381 30147 8415
rect 30147 8381 30156 8415
rect 30104 8372 30156 8381
rect 30196 8415 30248 8424
rect 30196 8381 30205 8415
rect 30205 8381 30239 8415
rect 30239 8381 30248 8415
rect 30196 8372 30248 8381
rect 31116 8372 31168 8424
rect 31392 8415 31444 8424
rect 31392 8381 31401 8415
rect 31401 8381 31435 8415
rect 31435 8381 31444 8415
rect 31392 8372 31444 8381
rect 31576 8415 31628 8424
rect 31576 8381 31585 8415
rect 31585 8381 31619 8415
rect 31619 8381 31628 8415
rect 31576 8372 31628 8381
rect 33232 8440 33284 8492
rect 33324 8415 33376 8424
rect 33324 8381 33333 8415
rect 33333 8381 33367 8415
rect 33367 8381 33376 8415
rect 33324 8372 33376 8381
rect 22928 8304 22980 8356
rect 24860 8347 24912 8356
rect 24860 8313 24878 8347
rect 24878 8313 24912 8347
rect 24860 8304 24912 8313
rect 29552 8304 29604 8356
rect 31484 8347 31536 8356
rect 31484 8313 31493 8347
rect 31493 8313 31527 8347
rect 31527 8313 31536 8347
rect 31484 8304 31536 8313
rect 32956 8304 33008 8356
rect 33140 8304 33192 8356
rect 23480 8279 23532 8288
rect 23480 8245 23489 8279
rect 23489 8245 23523 8279
rect 23523 8245 23532 8279
rect 23480 8236 23532 8245
rect 23756 8279 23808 8288
rect 23756 8245 23765 8279
rect 23765 8245 23799 8279
rect 23799 8245 23808 8279
rect 23756 8236 23808 8245
rect 12052 8134 12104 8186
rect 12116 8134 12168 8186
rect 12180 8134 12232 8186
rect 12244 8134 12296 8186
rect 23123 8134 23175 8186
rect 23187 8134 23239 8186
rect 23251 8134 23303 8186
rect 23315 8134 23367 8186
rect 3240 8032 3292 8084
rect 5356 8032 5408 8084
rect 5632 8032 5684 8084
rect 2320 7964 2372 8016
rect 1492 7896 1544 7948
rect 4528 7939 4580 7948
rect 4528 7905 4537 7939
rect 4537 7905 4571 7939
rect 4571 7905 4580 7939
rect 4528 7896 4580 7905
rect 8208 8032 8260 8084
rect 10416 8075 10468 8084
rect 10416 8041 10425 8075
rect 10425 8041 10459 8075
rect 10459 8041 10468 8075
rect 10416 8032 10468 8041
rect 10692 8032 10744 8084
rect 12992 8032 13044 8084
rect 13452 8075 13504 8084
rect 13452 8041 13461 8075
rect 13461 8041 13495 8075
rect 13495 8041 13504 8075
rect 13452 8032 13504 8041
rect 16120 8075 16172 8084
rect 16120 8041 16129 8075
rect 16129 8041 16163 8075
rect 16163 8041 16172 8075
rect 16120 8032 16172 8041
rect 17408 8032 17460 8084
rect 18328 8032 18380 8084
rect 24860 8032 24912 8084
rect 28540 8032 28592 8084
rect 29920 8032 29972 8084
rect 33140 8032 33192 8084
rect 9312 7964 9364 8016
rect 10784 8007 10836 8016
rect 8576 7896 8628 7948
rect 9956 7939 10008 7948
rect 9956 7905 9965 7939
rect 9965 7905 9999 7939
rect 9999 7905 10008 7939
rect 9956 7896 10008 7905
rect 10784 7973 10793 8007
rect 10793 7973 10827 8007
rect 10827 7973 10836 8007
rect 10784 7964 10836 7973
rect 2780 7828 2832 7880
rect 5172 7828 5224 7880
rect 8852 7828 8904 7880
rect 9588 7828 9640 7880
rect 12624 7896 12676 7948
rect 12900 7896 12952 7948
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 13544 7871 13596 7880
rect 10140 7760 10192 7812
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 15476 7896 15528 7948
rect 14740 7871 14792 7880
rect 14740 7837 14749 7871
rect 14749 7837 14783 7871
rect 14783 7837 14792 7871
rect 14740 7828 14792 7837
rect 18052 7896 18104 7948
rect 20352 7896 20404 7948
rect 21640 7939 21692 7948
rect 21640 7905 21674 7939
rect 21674 7905 21692 7939
rect 21640 7896 21692 7905
rect 23756 7896 23808 7948
rect 26976 7896 27028 7948
rect 27804 7939 27856 7948
rect 27804 7905 27813 7939
rect 27813 7905 27847 7939
rect 27847 7905 27856 7939
rect 27804 7896 27856 7905
rect 28172 7896 28224 7948
rect 29000 7964 29052 8016
rect 29552 8007 29604 8016
rect 29552 7973 29561 8007
rect 29561 7973 29595 8007
rect 29595 7973 29604 8007
rect 29552 7964 29604 7973
rect 29644 7964 29696 8016
rect 29276 7939 29328 7948
rect 29276 7905 29285 7939
rect 29285 7905 29319 7939
rect 29319 7905 29328 7939
rect 29276 7896 29328 7905
rect 30012 7896 30064 7948
rect 31116 7896 31168 7948
rect 31300 7939 31352 7948
rect 31300 7905 31309 7939
rect 31309 7905 31343 7939
rect 31343 7905 31352 7939
rect 31300 7896 31352 7905
rect 32312 7939 32364 7948
rect 32312 7905 32321 7939
rect 32321 7905 32355 7939
rect 32355 7905 32364 7939
rect 32312 7896 32364 7905
rect 33416 7896 33468 7948
rect 33600 7939 33652 7948
rect 33600 7905 33609 7939
rect 33609 7905 33643 7939
rect 33643 7905 33652 7939
rect 33600 7896 33652 7905
rect 16580 7760 16632 7812
rect 17960 7828 18012 7880
rect 21088 7828 21140 7880
rect 24124 7871 24176 7880
rect 24124 7837 24133 7871
rect 24133 7837 24167 7871
rect 24167 7837 24176 7871
rect 24124 7828 24176 7837
rect 29920 7828 29972 7880
rect 31208 7828 31260 7880
rect 31576 7828 31628 7880
rect 32404 7871 32456 7880
rect 32404 7837 32413 7871
rect 32413 7837 32447 7871
rect 32447 7837 32456 7871
rect 32404 7828 32456 7837
rect 7564 7692 7616 7744
rect 9772 7735 9824 7744
rect 9772 7701 9781 7735
rect 9781 7701 9815 7735
rect 9815 7701 9824 7735
rect 9772 7692 9824 7701
rect 11980 7735 12032 7744
rect 11980 7701 11989 7735
rect 11989 7701 12023 7735
rect 12023 7701 12032 7735
rect 11980 7692 12032 7701
rect 16672 7735 16724 7744
rect 16672 7701 16681 7735
rect 16681 7701 16715 7735
rect 16715 7701 16724 7735
rect 16672 7692 16724 7701
rect 17316 7692 17368 7744
rect 19616 7692 19668 7744
rect 23848 7760 23900 7812
rect 30104 7760 30156 7812
rect 22376 7692 22428 7744
rect 22468 7692 22520 7744
rect 33232 7692 33284 7744
rect 6517 7590 6569 7642
rect 6581 7590 6633 7642
rect 6645 7590 6697 7642
rect 6709 7590 6761 7642
rect 17588 7590 17640 7642
rect 17652 7590 17704 7642
rect 17716 7590 17768 7642
rect 17780 7590 17832 7642
rect 28658 7590 28710 7642
rect 28722 7590 28774 7642
rect 28786 7590 28838 7642
rect 28850 7590 28902 7642
rect 5172 7531 5224 7540
rect 5172 7497 5181 7531
rect 5181 7497 5215 7531
rect 5215 7497 5224 7531
rect 5172 7488 5224 7497
rect 8576 7488 8628 7540
rect 8668 7488 8720 7540
rect 15476 7488 15528 7540
rect 19708 7531 19760 7540
rect 19708 7497 19717 7531
rect 19717 7497 19751 7531
rect 19751 7497 19760 7531
rect 19708 7488 19760 7497
rect 21180 7488 21232 7540
rect 21640 7488 21692 7540
rect 23572 7488 23624 7540
rect 24124 7531 24176 7540
rect 24124 7497 24133 7531
rect 24133 7497 24167 7531
rect 24167 7497 24176 7531
rect 24124 7488 24176 7497
rect 4436 7420 4488 7472
rect 5448 7420 5500 7472
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 3332 7352 3384 7404
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 5632 7352 5684 7361
rect 22376 7420 22428 7472
rect 8300 7352 8352 7404
rect 10232 7395 10284 7404
rect 2964 7284 3016 7336
rect 7564 7327 7616 7336
rect 7564 7293 7573 7327
rect 7573 7293 7607 7327
rect 7607 7293 7616 7327
rect 7564 7284 7616 7293
rect 9036 7327 9088 7336
rect 9036 7293 9045 7327
rect 9045 7293 9079 7327
rect 9079 7293 9088 7327
rect 9036 7284 9088 7293
rect 9404 7284 9456 7336
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 9772 7284 9824 7336
rect 13452 7352 13504 7404
rect 15568 7395 15620 7404
rect 10784 7284 10836 7336
rect 11980 7284 12032 7336
rect 13268 7284 13320 7336
rect 13820 7327 13872 7336
rect 13820 7293 13829 7327
rect 13829 7293 13863 7327
rect 13863 7293 13872 7327
rect 13820 7284 13872 7293
rect 15568 7361 15577 7395
rect 15577 7361 15611 7395
rect 15611 7361 15620 7395
rect 15568 7352 15620 7361
rect 15752 7327 15804 7336
rect 15752 7293 15761 7327
rect 15761 7293 15795 7327
rect 15795 7293 15804 7327
rect 15752 7284 15804 7293
rect 16672 7284 16724 7336
rect 17132 7284 17184 7336
rect 17408 7284 17460 7336
rect 19616 7327 19668 7336
rect 19616 7293 19625 7327
rect 19625 7293 19659 7327
rect 19659 7293 19668 7327
rect 19616 7284 19668 7293
rect 19800 7327 19852 7336
rect 19800 7293 19809 7327
rect 19809 7293 19843 7327
rect 19843 7293 19852 7327
rect 19800 7284 19852 7293
rect 21364 7327 21416 7336
rect 21364 7293 21373 7327
rect 21373 7293 21407 7327
rect 21407 7293 21416 7327
rect 21364 7284 21416 7293
rect 22284 7284 22336 7336
rect 12716 7216 12768 7268
rect 1860 7148 1912 7200
rect 3240 7148 3292 7200
rect 5540 7191 5592 7200
rect 5540 7157 5549 7191
rect 5549 7157 5583 7191
rect 5583 7157 5592 7191
rect 5540 7148 5592 7157
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 9588 7148 9640 7200
rect 11796 7148 11848 7200
rect 14004 7191 14056 7200
rect 14004 7157 14013 7191
rect 14013 7157 14047 7191
rect 14047 7157 14056 7191
rect 14004 7148 14056 7157
rect 18052 7148 18104 7200
rect 22468 7216 22520 7268
rect 22928 7284 22980 7336
rect 25872 7420 25924 7472
rect 23480 7352 23532 7404
rect 23756 7284 23808 7336
rect 22928 7148 22980 7200
rect 28080 7284 28132 7336
rect 29920 7531 29972 7540
rect 29920 7497 29929 7531
rect 29929 7497 29963 7531
rect 29963 7497 29972 7531
rect 29920 7488 29972 7497
rect 32404 7488 32456 7540
rect 28540 7420 28592 7472
rect 29828 7420 29880 7472
rect 30012 7420 30064 7472
rect 33416 7463 33468 7472
rect 33416 7429 33425 7463
rect 33425 7429 33459 7463
rect 33459 7429 33468 7463
rect 33416 7420 33468 7429
rect 30472 7352 30524 7404
rect 31116 7352 31168 7404
rect 28448 7284 28500 7336
rect 29092 7327 29144 7336
rect 29092 7293 29101 7327
rect 29101 7293 29135 7327
rect 29135 7293 29144 7327
rect 29092 7284 29144 7293
rect 29552 7284 29604 7336
rect 30564 7327 30616 7336
rect 28724 7259 28776 7268
rect 28724 7225 28733 7259
rect 28733 7225 28767 7259
rect 28767 7225 28776 7259
rect 28724 7216 28776 7225
rect 29736 7216 29788 7268
rect 30564 7293 30573 7327
rect 30573 7293 30607 7327
rect 30607 7293 30616 7327
rect 30564 7284 30616 7293
rect 31208 7327 31260 7336
rect 31208 7293 31217 7327
rect 31217 7293 31251 7327
rect 31251 7293 31260 7327
rect 31208 7284 31260 7293
rect 31300 7327 31352 7336
rect 31300 7293 31309 7327
rect 31309 7293 31343 7327
rect 31343 7293 31352 7327
rect 31300 7284 31352 7293
rect 26056 7148 26108 7200
rect 26240 7148 26292 7200
rect 31392 7148 31444 7200
rect 33324 7216 33376 7268
rect 12052 7046 12104 7098
rect 12116 7046 12168 7098
rect 12180 7046 12232 7098
rect 12244 7046 12296 7098
rect 23123 7046 23175 7098
rect 23187 7046 23239 7098
rect 23251 7046 23303 7098
rect 23315 7046 23367 7098
rect 2320 6944 2372 6996
rect 2688 6944 2740 6996
rect 10784 6944 10836 6996
rect 13544 6944 13596 6996
rect 17960 6944 18012 6996
rect 28724 6944 28776 6996
rect 33600 6987 33652 6996
rect 33600 6953 33609 6987
rect 33609 6953 33643 6987
rect 33643 6953 33652 6987
rect 33600 6944 33652 6953
rect 5632 6876 5684 6928
rect 10600 6876 10652 6928
rect 13268 6876 13320 6928
rect 17132 6876 17184 6928
rect 18696 6876 18748 6928
rect 19524 6876 19576 6928
rect 1860 6851 1912 6860
rect 1860 6817 1869 6851
rect 1869 6817 1903 6851
rect 1903 6817 1912 6851
rect 1860 6808 1912 6817
rect 5540 6808 5592 6860
rect 11336 6808 11388 6860
rect 12716 6851 12768 6860
rect 12716 6817 12725 6851
rect 12725 6817 12759 6851
rect 12759 6817 12768 6851
rect 12716 6808 12768 6817
rect 1400 6740 1452 6792
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 10968 6740 11020 6792
rect 4528 6672 4580 6724
rect 10048 6672 10100 6724
rect 11612 6740 11664 6792
rect 13176 6808 13228 6860
rect 13636 6808 13688 6860
rect 15936 6808 15988 6860
rect 16212 6808 16264 6860
rect 16764 6851 16816 6860
rect 16764 6817 16773 6851
rect 16773 6817 16807 6851
rect 16807 6817 16816 6851
rect 16764 6808 16816 6817
rect 16488 6740 16540 6792
rect 13360 6672 13412 6724
rect 13544 6672 13596 6724
rect 15384 6672 15436 6724
rect 18052 6851 18104 6860
rect 18052 6817 18061 6851
rect 18061 6817 18095 6851
rect 18095 6817 18104 6851
rect 18052 6808 18104 6817
rect 19064 6851 19116 6860
rect 19064 6817 19073 6851
rect 19073 6817 19107 6851
rect 19107 6817 19116 6851
rect 19064 6808 19116 6817
rect 21272 6851 21324 6860
rect 21272 6817 21281 6851
rect 21281 6817 21315 6851
rect 21315 6817 21324 6851
rect 21272 6808 21324 6817
rect 23480 6808 23532 6860
rect 23940 6808 23992 6860
rect 25964 6876 26016 6928
rect 32588 6876 32640 6928
rect 26976 6808 27028 6860
rect 27804 6851 27856 6860
rect 20076 6740 20128 6792
rect 20352 6783 20404 6792
rect 20352 6749 20361 6783
rect 20361 6749 20395 6783
rect 20395 6749 20404 6783
rect 20352 6740 20404 6749
rect 23848 6783 23900 6792
rect 23848 6749 23857 6783
rect 23857 6749 23891 6783
rect 23891 6749 23900 6783
rect 23848 6740 23900 6749
rect 24032 6783 24084 6792
rect 24032 6749 24041 6783
rect 24041 6749 24075 6783
rect 24075 6749 24084 6783
rect 24032 6740 24084 6749
rect 26240 6740 26292 6792
rect 27804 6817 27813 6851
rect 27813 6817 27847 6851
rect 27847 6817 27856 6851
rect 27804 6808 27856 6817
rect 29276 6808 29328 6860
rect 29368 6851 29420 6860
rect 29368 6817 29377 6851
rect 29377 6817 29411 6851
rect 29411 6817 29420 6851
rect 29368 6808 29420 6817
rect 30012 6808 30064 6860
rect 31024 6740 31076 6792
rect 31576 6740 31628 6792
rect 33140 6740 33192 6792
rect 19616 6672 19668 6724
rect 2964 6604 3016 6656
rect 4252 6604 4304 6656
rect 12348 6604 12400 6656
rect 15568 6647 15620 6656
rect 15568 6613 15577 6647
rect 15577 6613 15611 6647
rect 15611 6613 15620 6647
rect 15568 6604 15620 6613
rect 15752 6604 15804 6656
rect 18696 6604 18748 6656
rect 18880 6647 18932 6656
rect 18880 6613 18889 6647
rect 18889 6613 18923 6647
rect 18923 6613 18932 6647
rect 18880 6604 18932 6613
rect 18972 6647 19024 6656
rect 18972 6613 18981 6647
rect 18981 6613 19015 6647
rect 19015 6613 19024 6647
rect 22560 6672 22612 6724
rect 18972 6604 19024 6613
rect 20260 6604 20312 6656
rect 21732 6647 21784 6656
rect 21732 6613 21741 6647
rect 21741 6613 21775 6647
rect 21775 6613 21784 6647
rect 21732 6604 21784 6613
rect 24400 6604 24452 6656
rect 28264 6604 28316 6656
rect 6517 6502 6569 6554
rect 6581 6502 6633 6554
rect 6645 6502 6697 6554
rect 6709 6502 6761 6554
rect 17588 6502 17640 6554
rect 17652 6502 17704 6554
rect 17716 6502 17768 6554
rect 17780 6502 17832 6554
rect 28658 6502 28710 6554
rect 28722 6502 28774 6554
rect 28786 6502 28838 6554
rect 28850 6502 28902 6554
rect 5540 6400 5592 6452
rect 9404 6443 9456 6452
rect 9404 6409 9413 6443
rect 9413 6409 9447 6443
rect 9447 6409 9456 6443
rect 9404 6400 9456 6409
rect 10968 6443 11020 6452
rect 10968 6409 10977 6443
rect 10977 6409 11011 6443
rect 11011 6409 11020 6443
rect 10968 6400 11020 6409
rect 4252 6307 4304 6316
rect 4252 6273 4261 6307
rect 4261 6273 4295 6307
rect 4295 6273 4304 6307
rect 4252 6264 4304 6273
rect 4528 6264 4580 6316
rect 6920 6307 6972 6316
rect 6920 6273 6929 6307
rect 6929 6273 6963 6307
rect 6963 6273 6972 6307
rect 6920 6264 6972 6273
rect 7196 6307 7248 6316
rect 7196 6273 7205 6307
rect 7205 6273 7239 6307
rect 7239 6273 7248 6307
rect 7196 6264 7248 6273
rect 10048 6307 10100 6316
rect 10048 6273 10057 6307
rect 10057 6273 10091 6307
rect 10091 6273 10100 6307
rect 10048 6264 10100 6273
rect 13176 6400 13228 6452
rect 13452 6400 13504 6452
rect 13544 6400 13596 6452
rect 16212 6443 16264 6452
rect 12808 6375 12860 6384
rect 12808 6341 12817 6375
rect 12817 6341 12851 6375
rect 12851 6341 12860 6375
rect 12808 6332 12860 6341
rect 13728 6332 13780 6384
rect 8208 6196 8260 6248
rect 5264 6128 5316 6180
rect 9496 6128 9548 6180
rect 10232 6196 10284 6248
rect 12624 6196 12676 6248
rect 13636 6264 13688 6316
rect 16212 6409 16221 6443
rect 16221 6409 16255 6443
rect 16255 6409 16264 6443
rect 16212 6400 16264 6409
rect 14740 6264 14792 6316
rect 19524 6307 19576 6316
rect 19524 6273 19533 6307
rect 19533 6273 19567 6307
rect 19567 6273 19576 6307
rect 21088 6400 21140 6452
rect 21732 6400 21784 6452
rect 22560 6400 22612 6452
rect 29276 6443 29328 6452
rect 29276 6409 29285 6443
rect 29285 6409 29319 6443
rect 29319 6409 29328 6443
rect 29276 6400 29328 6409
rect 29368 6400 29420 6452
rect 30564 6400 30616 6452
rect 33140 6400 33192 6452
rect 19524 6264 19576 6273
rect 23020 6264 23072 6316
rect 23664 6264 23716 6316
rect 14004 6196 14056 6248
rect 15568 6196 15620 6248
rect 18880 6196 18932 6248
rect 20260 6239 20312 6248
rect 20260 6205 20294 6239
rect 20294 6205 20312 6239
rect 20260 6196 20312 6205
rect 29276 6264 29328 6316
rect 13084 6128 13136 6180
rect 16120 6128 16172 6180
rect 22468 6128 22520 6180
rect 24400 6196 24452 6248
rect 28080 6239 28132 6248
rect 28080 6205 28089 6239
rect 28089 6205 28123 6239
rect 28123 6205 28132 6239
rect 28080 6196 28132 6205
rect 28264 6239 28316 6248
rect 28264 6205 28273 6239
rect 28273 6205 28307 6239
rect 28307 6205 28316 6239
rect 28264 6196 28316 6205
rect 28448 6196 28500 6248
rect 26056 6128 26108 6180
rect 30472 6196 30524 6248
rect 31668 6196 31720 6248
rect 32956 6196 33008 6248
rect 33232 6239 33284 6248
rect 33232 6205 33241 6239
rect 33241 6205 33275 6239
rect 33275 6205 33284 6239
rect 33232 6196 33284 6205
rect 29644 6128 29696 6180
rect 29736 6128 29788 6180
rect 9772 6103 9824 6112
rect 9772 6069 9781 6103
rect 9781 6069 9815 6103
rect 9815 6069 9824 6103
rect 9772 6060 9824 6069
rect 18420 6060 18472 6112
rect 21364 6103 21416 6112
rect 21364 6069 21373 6103
rect 21373 6069 21407 6103
rect 21407 6069 21416 6103
rect 21364 6060 21416 6069
rect 22560 6103 22612 6112
rect 22560 6069 22569 6103
rect 22569 6069 22603 6103
rect 22603 6069 22612 6103
rect 22560 6060 22612 6069
rect 25964 6060 26016 6112
rect 27804 6060 27856 6112
rect 31300 6128 31352 6180
rect 31668 6060 31720 6112
rect 12052 5958 12104 6010
rect 12116 5958 12168 6010
rect 12180 5958 12232 6010
rect 12244 5958 12296 6010
rect 23123 5958 23175 6010
rect 23187 5958 23239 6010
rect 23251 5958 23303 6010
rect 23315 5958 23367 6010
rect 2964 5899 3016 5908
rect 2964 5865 2973 5899
rect 2973 5865 3007 5899
rect 3007 5865 3016 5899
rect 2964 5856 3016 5865
rect 5632 5856 5684 5908
rect 9772 5856 9824 5908
rect 5264 5788 5316 5840
rect 12624 5856 12676 5908
rect 15936 5899 15988 5908
rect 15936 5865 15945 5899
rect 15945 5865 15979 5899
rect 15979 5865 15988 5899
rect 15936 5856 15988 5865
rect 16488 5899 16540 5908
rect 16488 5865 16497 5899
rect 16497 5865 16531 5899
rect 16531 5865 16540 5899
rect 16488 5856 16540 5865
rect 20076 5899 20128 5908
rect 20076 5865 20085 5899
rect 20085 5865 20119 5899
rect 20119 5865 20128 5899
rect 20076 5856 20128 5865
rect 20352 5856 20404 5908
rect 11796 5831 11848 5840
rect 11796 5797 11805 5831
rect 11805 5797 11839 5831
rect 11839 5797 11848 5831
rect 11796 5788 11848 5797
rect 13084 5788 13136 5840
rect 13728 5788 13780 5840
rect 16212 5788 16264 5840
rect 8576 5763 8628 5772
rect 8576 5729 8585 5763
rect 8585 5729 8619 5763
rect 8619 5729 8628 5763
rect 8576 5720 8628 5729
rect 9496 5720 9548 5772
rect 10232 5720 10284 5772
rect 10416 5763 10468 5772
rect 10416 5729 10425 5763
rect 10425 5729 10459 5763
rect 10459 5729 10468 5763
rect 10416 5720 10468 5729
rect 16120 5720 16172 5772
rect 22192 5788 22244 5840
rect 22560 5788 22612 5840
rect 26976 5856 27028 5908
rect 27528 5856 27580 5908
rect 29276 5899 29328 5908
rect 27804 5831 27856 5840
rect 27804 5797 27813 5831
rect 27813 5797 27847 5831
rect 27847 5797 27856 5831
rect 27804 5788 27856 5797
rect 29276 5865 29285 5899
rect 29285 5865 29319 5899
rect 29319 5865 29328 5899
rect 29276 5856 29328 5865
rect 30380 5788 30432 5840
rect 31484 5788 31536 5840
rect 32864 5788 32916 5840
rect 3056 5695 3108 5704
rect 3056 5661 3065 5695
rect 3065 5661 3099 5695
rect 3099 5661 3108 5695
rect 3056 5652 3108 5661
rect 3240 5695 3292 5704
rect 3240 5661 3249 5695
rect 3249 5661 3283 5695
rect 3283 5661 3292 5695
rect 3240 5652 3292 5661
rect 7104 5695 7156 5704
rect 7104 5661 7113 5695
rect 7113 5661 7147 5695
rect 7147 5661 7156 5695
rect 7104 5652 7156 5661
rect 9312 5652 9364 5704
rect 12348 5652 12400 5704
rect 14740 5652 14792 5704
rect 15384 5652 15436 5704
rect 17408 5763 17460 5772
rect 17408 5729 17417 5763
rect 17417 5729 17451 5763
rect 17451 5729 17460 5763
rect 17408 5720 17460 5729
rect 17960 5720 18012 5772
rect 18420 5720 18472 5772
rect 19616 5652 19668 5704
rect 21364 5720 21416 5772
rect 24308 5720 24360 5772
rect 25596 5695 25648 5704
rect 17316 5584 17368 5636
rect 17500 5627 17552 5636
rect 17500 5593 17509 5627
rect 17509 5593 17543 5627
rect 17543 5593 17552 5627
rect 17500 5584 17552 5593
rect 21732 5584 21784 5636
rect 2596 5559 2648 5568
rect 2596 5525 2605 5559
rect 2605 5525 2639 5559
rect 2639 5525 2648 5559
rect 2596 5516 2648 5525
rect 13360 5516 13412 5568
rect 18144 5559 18196 5568
rect 18144 5525 18153 5559
rect 18153 5525 18187 5559
rect 18187 5525 18196 5559
rect 18144 5516 18196 5525
rect 19064 5516 19116 5568
rect 23480 5559 23532 5568
rect 23480 5525 23489 5559
rect 23489 5525 23523 5559
rect 23523 5525 23532 5559
rect 23480 5516 23532 5525
rect 25596 5661 25605 5695
rect 25605 5661 25639 5695
rect 25639 5661 25648 5695
rect 25596 5652 25648 5661
rect 26056 5652 26108 5704
rect 31576 5652 31628 5704
rect 32128 5695 32180 5704
rect 32128 5661 32137 5695
rect 32137 5661 32171 5695
rect 32171 5661 32180 5695
rect 32128 5652 32180 5661
rect 26056 5516 26108 5568
rect 27068 5559 27120 5568
rect 27068 5525 27077 5559
rect 27077 5525 27111 5559
rect 27111 5525 27120 5559
rect 27068 5516 27120 5525
rect 29092 5516 29144 5568
rect 32312 5516 32364 5568
rect 6517 5414 6569 5466
rect 6581 5414 6633 5466
rect 6645 5414 6697 5466
rect 6709 5414 6761 5466
rect 17588 5414 17640 5466
rect 17652 5414 17704 5466
rect 17716 5414 17768 5466
rect 17780 5414 17832 5466
rect 28658 5414 28710 5466
rect 28722 5414 28774 5466
rect 28786 5414 28838 5466
rect 28850 5414 28902 5466
rect 3056 5312 3108 5364
rect 7104 5312 7156 5364
rect 8576 5312 8628 5364
rect 10600 5355 10652 5364
rect 10600 5321 10609 5355
rect 10609 5321 10643 5355
rect 10643 5321 10652 5355
rect 10600 5312 10652 5321
rect 13636 5312 13688 5364
rect 20536 5312 20588 5364
rect 22192 5312 22244 5364
rect 23020 5312 23072 5364
rect 24032 5312 24084 5364
rect 25596 5312 25648 5364
rect 32128 5312 32180 5364
rect 25688 5244 25740 5296
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 2596 5176 2648 5228
rect 5356 5219 5408 5228
rect 5356 5185 5365 5219
rect 5365 5185 5399 5219
rect 5399 5185 5408 5219
rect 5356 5176 5408 5185
rect 5632 5176 5684 5228
rect 10324 5219 10376 5228
rect 10324 5185 10333 5219
rect 10333 5185 10367 5219
rect 10367 5185 10376 5219
rect 10324 5176 10376 5185
rect 16304 5176 16356 5228
rect 17132 5176 17184 5228
rect 20812 5176 20864 5228
rect 25964 5219 26016 5228
rect 2688 5108 2740 5160
rect 9404 5108 9456 5160
rect 5172 5040 5224 5092
rect 9220 5040 9272 5092
rect 10416 5108 10468 5160
rect 13360 5151 13412 5160
rect 13360 5117 13369 5151
rect 13369 5117 13403 5151
rect 13403 5117 13412 5151
rect 13360 5108 13412 5117
rect 17408 5108 17460 5160
rect 21364 5151 21416 5160
rect 16488 5040 16540 5092
rect 21364 5117 21373 5151
rect 21373 5117 21407 5151
rect 21407 5117 21416 5151
rect 21364 5108 21416 5117
rect 22928 5108 22980 5160
rect 23480 5108 23532 5160
rect 25964 5185 25973 5219
rect 25973 5185 26007 5219
rect 26007 5185 26016 5219
rect 25964 5176 26016 5185
rect 31300 5244 31352 5296
rect 24308 5151 24360 5160
rect 24308 5117 24317 5151
rect 24317 5117 24351 5151
rect 24351 5117 24360 5151
rect 24308 5108 24360 5117
rect 30380 5151 30432 5160
rect 30380 5117 30389 5151
rect 30389 5117 30423 5151
rect 30423 5117 30432 5151
rect 30380 5108 30432 5117
rect 32312 5176 32364 5228
rect 31668 5151 31720 5160
rect 31668 5117 31677 5151
rect 31677 5117 31711 5151
rect 31711 5117 31720 5151
rect 31668 5108 31720 5117
rect 31944 5151 31996 5160
rect 31944 5117 31953 5151
rect 31953 5117 31987 5151
rect 31987 5117 31996 5151
rect 31944 5108 31996 5117
rect 32956 5108 33008 5160
rect 33048 5108 33100 5160
rect 31484 5040 31536 5092
rect 5540 5015 5592 5024
rect 5540 4981 5549 5015
rect 5549 4981 5583 5015
rect 5583 4981 5592 5015
rect 5540 4972 5592 4981
rect 15016 4972 15068 5024
rect 16120 4972 16172 5024
rect 17960 4972 18012 5024
rect 20904 5015 20956 5024
rect 20904 4981 20913 5015
rect 20913 4981 20947 5015
rect 20947 4981 20956 5015
rect 20904 4972 20956 4981
rect 27068 4972 27120 5024
rect 30564 4972 30616 5024
rect 31852 4972 31904 5024
rect 33416 4972 33468 5024
rect 12052 4870 12104 4922
rect 12116 4870 12168 4922
rect 12180 4870 12232 4922
rect 12244 4870 12296 4922
rect 23123 4870 23175 4922
rect 23187 4870 23239 4922
rect 23251 4870 23303 4922
rect 23315 4870 23367 4922
rect 12992 4768 13044 4820
rect 13728 4768 13780 4820
rect 3056 4700 3108 4752
rect 5172 4700 5224 4752
rect 15016 4743 15068 4752
rect 15016 4709 15025 4743
rect 15025 4709 15059 4743
rect 15059 4709 15068 4743
rect 15016 4700 15068 4709
rect 17316 4768 17368 4820
rect 22376 4811 22428 4820
rect 22376 4777 22385 4811
rect 22385 4777 22419 4811
rect 22419 4777 22428 4811
rect 22376 4768 22428 4777
rect 31852 4768 31904 4820
rect 16304 4700 16356 4752
rect 4528 4632 4580 4684
rect 14740 4675 14792 4684
rect 14740 4641 14749 4675
rect 14749 4641 14783 4675
rect 14783 4641 14792 4675
rect 14740 4632 14792 4641
rect 17960 4675 18012 4684
rect 3056 4607 3108 4616
rect 3056 4573 3065 4607
rect 3065 4573 3099 4607
rect 3099 4573 3108 4607
rect 3056 4564 3108 4573
rect 3240 4607 3292 4616
rect 3240 4573 3249 4607
rect 3249 4573 3283 4607
rect 3283 4573 3292 4607
rect 3240 4564 3292 4573
rect 4620 4607 4672 4616
rect 4620 4573 4629 4607
rect 4629 4573 4663 4607
rect 4663 4573 4672 4607
rect 4620 4564 4672 4573
rect 17960 4641 17969 4675
rect 17969 4641 18003 4675
rect 18003 4641 18012 4675
rect 17960 4632 18012 4641
rect 18328 4632 18380 4684
rect 19156 4632 19208 4684
rect 19892 4632 19944 4684
rect 20168 4675 20220 4684
rect 20168 4641 20177 4675
rect 20177 4641 20211 4675
rect 20211 4641 20220 4675
rect 20168 4632 20220 4641
rect 20904 4700 20956 4752
rect 20720 4564 20772 4616
rect 24400 4632 24452 4684
rect 28080 4700 28132 4752
rect 28540 4700 28592 4752
rect 33416 4743 33468 4752
rect 27620 4675 27672 4684
rect 27620 4641 27629 4675
rect 27629 4641 27663 4675
rect 27663 4641 27672 4675
rect 27620 4632 27672 4641
rect 28448 4632 28500 4684
rect 30564 4675 30616 4684
rect 30564 4641 30573 4675
rect 30573 4641 30607 4675
rect 30607 4641 30616 4675
rect 30564 4632 30616 4641
rect 30748 4675 30800 4684
rect 30748 4641 30757 4675
rect 30757 4641 30791 4675
rect 30791 4641 30800 4675
rect 30748 4632 30800 4641
rect 31208 4675 31260 4684
rect 31208 4641 31217 4675
rect 31217 4641 31251 4675
rect 31251 4641 31260 4675
rect 31208 4632 31260 4641
rect 31852 4632 31904 4684
rect 33416 4709 33425 4743
rect 33425 4709 33459 4743
rect 33459 4709 33468 4743
rect 33416 4700 33468 4709
rect 33600 4743 33652 4752
rect 33600 4709 33609 4743
rect 33609 4709 33643 4743
rect 33643 4709 33652 4743
rect 33600 4700 33652 4709
rect 32312 4632 32364 4684
rect 25688 4564 25740 4616
rect 29460 4564 29512 4616
rect 33048 4564 33100 4616
rect 20628 4496 20680 4548
rect 27068 4496 27120 4548
rect 32496 4496 32548 4548
rect 1860 4471 1912 4480
rect 1860 4437 1869 4471
rect 1869 4437 1903 4471
rect 1903 4437 1912 4471
rect 1860 4428 1912 4437
rect 2596 4471 2648 4480
rect 2596 4437 2605 4471
rect 2605 4437 2639 4471
rect 2639 4437 2648 4471
rect 2596 4428 2648 4437
rect 5632 4428 5684 4480
rect 16488 4471 16540 4480
rect 16488 4437 16497 4471
rect 16497 4437 16531 4471
rect 16531 4437 16540 4471
rect 16488 4428 16540 4437
rect 18972 4471 19024 4480
rect 18972 4437 18981 4471
rect 18981 4437 19015 4471
rect 19015 4437 19024 4471
rect 18972 4428 19024 4437
rect 20996 4428 21048 4480
rect 22928 4428 22980 4480
rect 26792 4428 26844 4480
rect 31852 4428 31904 4480
rect 6517 4326 6569 4378
rect 6581 4326 6633 4378
rect 6645 4326 6697 4378
rect 6709 4326 6761 4378
rect 17588 4326 17640 4378
rect 17652 4326 17704 4378
rect 17716 4326 17768 4378
rect 17780 4326 17832 4378
rect 28658 4326 28710 4378
rect 28722 4326 28774 4378
rect 28786 4326 28838 4378
rect 28850 4326 28902 4378
rect 3056 4224 3108 4276
rect 4068 4224 4120 4276
rect 9588 4267 9640 4276
rect 9588 4233 9618 4267
rect 9618 4233 9640 4267
rect 9588 4224 9640 4233
rect 14648 4224 14700 4276
rect 20812 4224 20864 4276
rect 22928 4267 22980 4276
rect 22928 4233 22958 4267
rect 22958 4233 22980 4267
rect 22928 4224 22980 4233
rect 27620 4224 27672 4276
rect 28448 4224 28500 4276
rect 29460 4224 29512 4276
rect 31208 4224 31260 4276
rect 1400 4088 1452 4140
rect 2596 4088 2648 4140
rect 5356 4131 5408 4140
rect 5356 4097 5365 4131
rect 5365 4097 5399 4131
rect 5399 4097 5408 4131
rect 5356 4088 5408 4097
rect 5540 4088 5592 4140
rect 9312 4131 9364 4140
rect 9312 4097 9321 4131
rect 9321 4097 9355 4131
rect 9355 4097 9364 4131
rect 9312 4088 9364 4097
rect 10324 4088 10376 4140
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 14740 4131 14792 4140
rect 14740 4097 14749 4131
rect 14749 4097 14783 4131
rect 14783 4097 14792 4131
rect 14740 4088 14792 4097
rect 17132 4088 17184 4140
rect 18972 4020 19024 4072
rect 21088 4088 21140 4140
rect 22376 4088 22428 4140
rect 29092 4156 29144 4208
rect 20996 4063 21048 4072
rect 20996 4029 21005 4063
rect 21005 4029 21039 4063
rect 21039 4029 21048 4063
rect 20996 4020 21048 4029
rect 5172 3952 5224 4004
rect 5632 3952 5684 4004
rect 7012 3884 7064 3936
rect 13728 3952 13780 4004
rect 20720 3952 20772 4004
rect 27528 4020 27580 4072
rect 28540 4020 28592 4072
rect 28632 4020 28684 4072
rect 29460 4063 29512 4072
rect 29460 4029 29469 4063
rect 29469 4029 29503 4063
rect 29503 4029 29512 4063
rect 29460 4020 29512 4029
rect 30288 4063 30340 4072
rect 30288 4029 30297 4063
rect 30297 4029 30331 4063
rect 30331 4029 30340 4063
rect 30288 4020 30340 4029
rect 30748 4156 30800 4208
rect 31484 4131 31536 4140
rect 31484 4097 31493 4131
rect 31493 4097 31527 4131
rect 31527 4097 31536 4131
rect 31484 4088 31536 4097
rect 30748 4020 30800 4072
rect 31208 4063 31260 4072
rect 31208 4029 31217 4063
rect 31217 4029 31251 4063
rect 31251 4029 31260 4063
rect 31208 4020 31260 4029
rect 20168 3884 20220 3936
rect 28448 3952 28500 4004
rect 24400 3927 24452 3936
rect 24400 3893 24409 3927
rect 24409 3893 24443 3927
rect 24443 3893 24452 3927
rect 30380 3952 30432 4004
rect 24400 3884 24452 3893
rect 29092 3884 29144 3936
rect 29552 3884 29604 3936
rect 30196 3884 30248 3936
rect 12052 3782 12104 3834
rect 12116 3782 12168 3834
rect 12180 3782 12232 3834
rect 12244 3782 12296 3834
rect 23123 3782 23175 3834
rect 23187 3782 23239 3834
rect 23251 3782 23303 3834
rect 23315 3782 23367 3834
rect 4620 3680 4672 3732
rect 5540 3680 5592 3732
rect 6920 3680 6972 3732
rect 29552 3723 29604 3732
rect 5172 3612 5224 3664
rect 4068 3544 4120 3596
rect 5632 3544 5684 3596
rect 7012 3587 7064 3596
rect 7012 3553 7021 3587
rect 7021 3553 7055 3587
rect 7055 3553 7064 3587
rect 7012 3544 7064 3553
rect 29552 3689 29561 3723
rect 29561 3689 29595 3723
rect 29595 3689 29604 3723
rect 29552 3680 29604 3689
rect 31484 3680 31536 3732
rect 17132 3612 17184 3664
rect 26792 3655 26844 3664
rect 17408 3544 17460 3596
rect 26792 3621 26801 3655
rect 26801 3621 26835 3655
rect 26835 3621 26844 3655
rect 26792 3612 26844 3621
rect 27528 3612 27580 3664
rect 28540 3655 28592 3664
rect 28540 3621 28549 3655
rect 28549 3621 28583 3655
rect 28583 3621 28592 3655
rect 28540 3612 28592 3621
rect 18144 3587 18196 3596
rect 18144 3553 18153 3587
rect 18153 3553 18187 3587
rect 18187 3553 18196 3587
rect 18144 3544 18196 3553
rect 19156 3544 19208 3596
rect 21088 3544 21140 3596
rect 29184 3544 29236 3596
rect 31208 3612 31260 3664
rect 31852 3655 31904 3664
rect 31852 3621 31861 3655
rect 31861 3621 31895 3655
rect 31895 3621 31904 3655
rect 31852 3612 31904 3621
rect 32864 3612 32916 3664
rect 30748 3587 30800 3596
rect 5356 3476 5408 3528
rect 18420 3519 18472 3528
rect 18420 3485 18429 3519
rect 18429 3485 18463 3519
rect 18463 3485 18472 3519
rect 18420 3476 18472 3485
rect 26516 3519 26568 3528
rect 26516 3485 26525 3519
rect 26525 3485 26559 3519
rect 26559 3485 26568 3519
rect 26516 3476 26568 3485
rect 16120 3383 16172 3392
rect 16120 3349 16129 3383
rect 16129 3349 16163 3383
rect 16163 3349 16172 3383
rect 16120 3340 16172 3349
rect 18328 3383 18380 3392
rect 18328 3349 18337 3383
rect 18337 3349 18371 3383
rect 18371 3349 18380 3383
rect 18328 3340 18380 3349
rect 20444 3340 20496 3392
rect 30748 3553 30757 3587
rect 30757 3553 30791 3587
rect 30791 3553 30800 3587
rect 30748 3544 30800 3553
rect 31576 3587 31628 3596
rect 31576 3553 31585 3587
rect 31585 3553 31619 3587
rect 31619 3553 31628 3587
rect 31576 3544 31628 3553
rect 30288 3476 30340 3528
rect 30196 3340 30248 3392
rect 6517 3238 6569 3290
rect 6581 3238 6633 3290
rect 6645 3238 6697 3290
rect 6709 3238 6761 3290
rect 17588 3238 17640 3290
rect 17652 3238 17704 3290
rect 17716 3238 17768 3290
rect 17780 3238 17832 3290
rect 28658 3238 28710 3290
rect 28722 3238 28774 3290
rect 28786 3238 28838 3290
rect 28850 3238 28902 3290
rect 17408 3136 17460 3188
rect 19156 3136 19208 3188
rect 26516 3136 26568 3188
rect 17592 3043 17644 3052
rect 17592 3009 17601 3043
rect 17601 3009 17635 3043
rect 17635 3009 17644 3043
rect 17592 3000 17644 3009
rect 30288 3136 30340 3188
rect 31208 3136 31260 3188
rect 31576 3068 31628 3120
rect 29092 3000 29144 3052
rect 17224 2932 17276 2984
rect 18328 2975 18380 2984
rect 18328 2941 18362 2975
rect 18362 2941 18380 2975
rect 17132 2864 17184 2916
rect 18328 2932 18380 2941
rect 20444 2975 20496 2984
rect 20444 2941 20453 2975
rect 20453 2941 20487 2975
rect 20487 2941 20496 2975
rect 20444 2932 20496 2941
rect 19432 2839 19484 2848
rect 19432 2805 19441 2839
rect 19441 2805 19475 2839
rect 19475 2805 19484 2839
rect 19432 2796 19484 2805
rect 19892 2864 19944 2916
rect 21916 2932 21968 2984
rect 30656 2975 30708 2984
rect 30656 2941 30665 2975
rect 30665 2941 30699 2975
rect 30699 2941 30708 2975
rect 30656 2932 30708 2941
rect 20536 2796 20588 2848
rect 20720 2839 20772 2848
rect 20720 2805 20729 2839
rect 20729 2805 20763 2839
rect 20763 2805 20772 2839
rect 20720 2796 20772 2805
rect 27528 2796 27580 2848
rect 32864 2864 32916 2916
rect 12052 2694 12104 2746
rect 12116 2694 12168 2746
rect 12180 2694 12232 2746
rect 12244 2694 12296 2746
rect 23123 2694 23175 2746
rect 23187 2694 23239 2746
rect 23251 2694 23303 2746
rect 23315 2694 23367 2746
rect 5724 2635 5776 2644
rect 5724 2601 5733 2635
rect 5733 2601 5767 2635
rect 5767 2601 5776 2635
rect 5724 2592 5776 2601
rect 11244 2567 11296 2576
rect 11244 2533 11253 2567
rect 11253 2533 11287 2567
rect 11287 2533 11296 2567
rect 11244 2524 11296 2533
rect 12440 2592 12492 2644
rect 17592 2592 17644 2644
rect 18420 2635 18472 2644
rect 18420 2601 18429 2635
rect 18429 2601 18463 2635
rect 18463 2601 18472 2635
rect 18420 2592 18472 2601
rect 21916 2635 21968 2644
rect 21916 2601 21925 2635
rect 21925 2601 21959 2635
rect 21959 2601 21968 2635
rect 21916 2592 21968 2601
rect 16028 2524 16080 2576
rect 16488 2567 16540 2576
rect 16488 2533 16497 2567
rect 16497 2533 16531 2567
rect 16531 2533 16540 2567
rect 16488 2524 16540 2533
rect 2780 2456 2832 2508
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 13820 2456 13872 2508
rect 480 2320 532 2372
rect 16120 2388 16172 2440
rect 19432 2524 19484 2576
rect 20720 2524 20772 2576
rect 25780 2567 25832 2576
rect 25780 2533 25789 2567
rect 25789 2533 25823 2567
rect 25823 2533 25832 2567
rect 25780 2524 25832 2533
rect 28448 2567 28500 2576
rect 28448 2533 28457 2567
rect 28457 2533 28491 2567
rect 28491 2533 28500 2567
rect 28448 2524 28500 2533
rect 30380 2524 30432 2576
rect 31760 2567 31812 2576
rect 31760 2533 31769 2567
rect 31769 2533 31803 2567
rect 31803 2533 31812 2567
rect 31760 2524 31812 2533
rect 32496 2567 32548 2576
rect 32496 2533 32505 2567
rect 32505 2533 32539 2567
rect 32539 2533 32548 2567
rect 32496 2524 32548 2533
rect 20536 2499 20588 2508
rect 20536 2465 20545 2499
rect 20545 2465 20579 2499
rect 20579 2465 20588 2499
rect 20536 2456 20588 2465
rect 19984 2388 20036 2440
rect 8300 2363 8352 2372
rect 8300 2329 8309 2363
rect 8309 2329 8343 2363
rect 8343 2329 8352 2363
rect 8300 2320 8352 2329
rect 11060 2363 11112 2372
rect 11060 2329 11069 2363
rect 11069 2329 11103 2363
rect 11103 2329 11112 2363
rect 11060 2320 11112 2329
rect 19340 2363 19392 2372
rect 19340 2329 19349 2363
rect 19349 2329 19383 2363
rect 19383 2329 19392 2363
rect 19340 2320 19392 2329
rect 22100 2320 22152 2372
rect 24860 2320 24912 2372
rect 27620 2320 27672 2372
rect 30380 2320 30432 2372
rect 31944 2363 31996 2372
rect 31944 2329 31953 2363
rect 31953 2329 31987 2363
rect 31987 2329 31996 2363
rect 31944 2320 31996 2329
rect 32680 2363 32732 2372
rect 32680 2329 32689 2363
rect 32689 2329 32723 2363
rect 32723 2329 32732 2363
rect 32680 2320 32732 2329
rect 16304 2252 16356 2304
rect 16580 2295 16632 2304
rect 16580 2261 16589 2295
rect 16589 2261 16623 2295
rect 16623 2261 16632 2295
rect 16580 2252 16632 2261
rect 6517 2150 6569 2202
rect 6581 2150 6633 2202
rect 6645 2150 6697 2202
rect 6709 2150 6761 2202
rect 17588 2150 17640 2202
rect 17652 2150 17704 2202
rect 17716 2150 17768 2202
rect 17780 2150 17832 2202
rect 28658 2150 28710 2202
rect 28722 2150 28774 2202
rect 28786 2150 28838 2202
rect 28850 2150 28902 2202
<< metal2 >>
rect 2778 36853 2834 37653
rect 5078 36853 5134 37653
rect 7838 36853 7894 37653
rect 10598 36853 10654 37653
rect 13358 36853 13414 37653
rect 16118 36853 16174 37653
rect 18878 36853 18934 37653
rect 21638 36853 21694 37653
rect 24398 36853 24454 37653
rect 27158 36853 27214 37653
rect 29918 36853 29974 37653
rect 32678 36853 32734 37653
rect 34978 36853 35034 37653
rect 1398 36816 1454 36825
rect 1398 36751 1454 36760
rect 1412 35154 1440 36751
rect 2792 35154 2820 36853
rect 5092 35154 5120 36853
rect 7104 35488 7156 35494
rect 7104 35430 7156 35436
rect 7116 35290 7144 35430
rect 7104 35284 7156 35290
rect 7104 35226 7156 35232
rect 7852 35154 7880 36853
rect 10612 35222 10640 36853
rect 12026 35388 12322 35408
rect 12082 35386 12106 35388
rect 12162 35386 12186 35388
rect 12242 35386 12266 35388
rect 12104 35334 12106 35386
rect 12168 35334 12180 35386
rect 12242 35334 12244 35386
rect 12082 35332 12106 35334
rect 12162 35332 12186 35334
rect 12242 35332 12266 35334
rect 12026 35312 12322 35332
rect 12624 35284 12676 35290
rect 12624 35226 12676 35232
rect 10600 35216 10652 35222
rect 10600 35158 10652 35164
rect 1400 35148 1452 35154
rect 1400 35090 1452 35096
rect 2780 35148 2832 35154
rect 2780 35090 2832 35096
rect 5080 35148 5132 35154
rect 5080 35090 5132 35096
rect 7840 35148 7892 35154
rect 7840 35090 7892 35096
rect 8392 35148 8444 35154
rect 8392 35090 8444 35096
rect 8208 35012 8260 35018
rect 8208 34954 8260 34960
rect 2964 34944 3016 34950
rect 2964 34886 3016 34892
rect 2976 34678 3004 34886
rect 6491 34844 6787 34864
rect 6547 34842 6571 34844
rect 6627 34842 6651 34844
rect 6707 34842 6731 34844
rect 6569 34790 6571 34842
rect 6633 34790 6645 34842
rect 6707 34790 6709 34842
rect 6547 34788 6571 34790
rect 6627 34788 6651 34790
rect 6707 34788 6731 34790
rect 6491 34768 6787 34788
rect 2964 34672 3016 34678
rect 2964 34614 3016 34620
rect 7196 34604 7248 34610
rect 7196 34546 7248 34552
rect 6491 33756 6787 33776
rect 6547 33754 6571 33756
rect 6627 33754 6651 33756
rect 6707 33754 6731 33756
rect 6569 33702 6571 33754
rect 6633 33702 6645 33754
rect 6707 33702 6709 33754
rect 6547 33700 6571 33702
rect 6627 33700 6651 33702
rect 6707 33700 6731 33702
rect 6491 33680 6787 33700
rect 5080 33516 5132 33522
rect 5080 33458 5132 33464
rect 2964 33448 3016 33454
rect 2964 33390 3016 33396
rect 3976 33448 4028 33454
rect 3976 33390 4028 33396
rect 1400 32972 1452 32978
rect 1400 32914 1452 32920
rect 1412 32745 1440 32914
rect 1398 32736 1454 32745
rect 1398 32671 1454 32680
rect 2976 30734 3004 33390
rect 3056 33380 3108 33386
rect 3056 33322 3108 33328
rect 3068 30734 3096 33322
rect 3608 33312 3660 33318
rect 3608 33254 3660 33260
rect 3620 32366 3648 33254
rect 3884 33040 3936 33046
rect 3884 32982 3936 32988
rect 3896 32366 3924 32982
rect 3608 32360 3660 32366
rect 3608 32302 3660 32308
rect 3884 32360 3936 32366
rect 3884 32302 3936 32308
rect 3148 32224 3200 32230
rect 3148 32166 3200 32172
rect 3160 31890 3188 32166
rect 3896 31958 3924 32302
rect 3988 32026 4016 33390
rect 4528 32768 4580 32774
rect 4528 32710 4580 32716
rect 4540 32230 4568 32710
rect 5092 32570 5120 33458
rect 5448 33380 5500 33386
rect 5448 33322 5500 33328
rect 5080 32564 5132 32570
rect 5080 32506 5132 32512
rect 5356 32428 5408 32434
rect 5356 32370 5408 32376
rect 4528 32224 4580 32230
rect 4528 32166 4580 32172
rect 3976 32020 4028 32026
rect 3976 31962 4028 31968
rect 3884 31952 3936 31958
rect 3884 31894 3936 31900
rect 3148 31884 3200 31890
rect 3148 31826 3200 31832
rect 3160 31346 3188 31826
rect 3148 31340 3200 31346
rect 3148 31282 3200 31288
rect 3700 31340 3752 31346
rect 3700 31282 3752 31288
rect 3148 31136 3200 31142
rect 3148 31078 3200 31084
rect 3160 30802 3188 31078
rect 3148 30796 3200 30802
rect 3148 30738 3200 30744
rect 2964 30728 3016 30734
rect 2964 30670 3016 30676
rect 3056 30728 3108 30734
rect 3056 30670 3108 30676
rect 3240 30728 3292 30734
rect 3240 30670 3292 30676
rect 2780 30592 2832 30598
rect 2780 30534 2832 30540
rect 2792 30190 2820 30534
rect 1400 30184 1452 30190
rect 1400 30126 1452 30132
rect 2780 30184 2832 30190
rect 2780 30126 2832 30132
rect 1412 28626 1440 30126
rect 3068 29102 3096 30670
rect 3148 30048 3200 30054
rect 3148 29990 3200 29996
rect 3160 29714 3188 29990
rect 3252 29850 3280 30670
rect 3712 30190 3740 31282
rect 3700 30184 3752 30190
rect 3700 30126 3752 30132
rect 3240 29844 3292 29850
rect 3240 29786 3292 29792
rect 3148 29708 3200 29714
rect 3148 29650 3200 29656
rect 3424 29504 3476 29510
rect 3424 29446 3476 29452
rect 3436 29170 3464 29446
rect 3240 29164 3292 29170
rect 3240 29106 3292 29112
rect 3424 29164 3476 29170
rect 3424 29106 3476 29112
rect 1768 29096 1820 29102
rect 1768 29038 1820 29044
rect 3056 29096 3108 29102
rect 3056 29038 3108 29044
rect 1780 28665 1808 29038
rect 3056 28960 3108 28966
rect 3056 28902 3108 28908
rect 3068 28694 3096 28902
rect 3056 28688 3108 28694
rect 1766 28656 1822 28665
rect 1400 28620 1452 28626
rect 3056 28630 3108 28636
rect 1766 28591 1822 28600
rect 1400 28562 1452 28568
rect 2964 27940 3016 27946
rect 2964 27882 3016 27888
rect 2976 27538 3004 27882
rect 2964 27532 3016 27538
rect 2964 27474 3016 27480
rect 2780 27464 2832 27470
rect 2780 27406 2832 27412
rect 2688 27328 2740 27334
rect 2688 27270 2740 27276
rect 1492 26988 1544 26994
rect 1492 26930 1544 26936
rect 1504 24750 1532 26930
rect 2700 26926 2728 27270
rect 2688 26920 2740 26926
rect 2688 26862 2740 26868
rect 1584 26512 1636 26518
rect 1584 26454 1636 26460
rect 1492 24744 1544 24750
rect 1492 24686 1544 24692
rect 1398 24576 1454 24585
rect 1398 24511 1454 24520
rect 1412 24274 1440 24511
rect 1400 24268 1452 24274
rect 1400 24210 1452 24216
rect 1504 24154 1532 24686
rect 1412 24126 1532 24154
rect 1412 23118 1440 24126
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1412 21486 1440 23054
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 1412 19310 1440 21422
rect 1400 19304 1452 19310
rect 1400 19246 1452 19252
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1412 14958 1440 15982
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1412 12782 1440 14894
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1412 11218 1440 12718
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 8265 1440 8366
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1504 7954 1532 9454
rect 1596 8634 1624 26454
rect 2792 25770 2820 27406
rect 2872 26784 2924 26790
rect 2872 26726 2924 26732
rect 2884 26450 2912 26726
rect 2872 26444 2924 26450
rect 2872 26386 2924 26392
rect 2780 25764 2832 25770
rect 2780 25706 2832 25712
rect 1768 25356 1820 25362
rect 1768 25298 1820 25304
rect 1780 24070 1808 25298
rect 2792 25294 2820 25706
rect 2976 25430 3004 27474
rect 3148 27464 3200 27470
rect 3148 27406 3200 27412
rect 3160 26586 3188 27406
rect 3148 26580 3200 26586
rect 3148 26522 3200 26528
rect 3252 25906 3280 29106
rect 3332 29096 3384 29102
rect 3332 29038 3384 29044
rect 3344 28218 3372 29038
rect 3896 28626 3924 31894
rect 4540 31890 4568 32166
rect 4528 31884 4580 31890
rect 4528 31826 4580 31832
rect 4344 31816 4396 31822
rect 4344 31758 4396 31764
rect 4356 31414 4384 31758
rect 4344 31408 4396 31414
rect 4344 31350 4396 31356
rect 4068 30660 4120 30666
rect 4068 30602 4120 30608
rect 4080 29238 4108 30602
rect 4252 30184 4304 30190
rect 4252 30126 4304 30132
rect 4068 29232 4120 29238
rect 4068 29174 4120 29180
rect 4264 29102 4292 30126
rect 4356 29730 4384 31350
rect 5368 31346 5396 32370
rect 5460 31822 5488 33322
rect 6920 33312 6972 33318
rect 6920 33254 6972 33260
rect 5632 32972 5684 32978
rect 5632 32914 5684 32920
rect 5540 32224 5592 32230
rect 5540 32166 5592 32172
rect 5448 31816 5500 31822
rect 5448 31758 5500 31764
rect 4988 31340 5040 31346
rect 4988 31282 5040 31288
rect 5356 31340 5408 31346
rect 5356 31282 5408 31288
rect 4804 30796 4856 30802
rect 4804 30738 4856 30744
rect 4816 30394 4844 30738
rect 5000 30734 5028 31282
rect 5460 30870 5488 31758
rect 5552 31278 5580 32166
rect 5644 32026 5672 32914
rect 6932 32774 6960 33254
rect 6920 32768 6972 32774
rect 6920 32710 6972 32716
rect 6491 32668 6787 32688
rect 6547 32666 6571 32668
rect 6627 32666 6651 32668
rect 6707 32666 6731 32668
rect 6569 32614 6571 32666
rect 6633 32614 6645 32666
rect 6707 32614 6709 32666
rect 6547 32612 6571 32614
rect 6627 32612 6651 32614
rect 6707 32612 6731 32614
rect 6491 32592 6787 32612
rect 6932 32366 6960 32710
rect 6920 32360 6972 32366
rect 6920 32302 6972 32308
rect 5724 32224 5776 32230
rect 5724 32166 5776 32172
rect 5632 32020 5684 32026
rect 5632 31962 5684 31968
rect 5736 31890 5764 32166
rect 6828 31952 6880 31958
rect 6828 31894 6880 31900
rect 5724 31884 5776 31890
rect 5724 31826 5776 31832
rect 5724 31748 5776 31754
rect 5724 31690 5776 31696
rect 5540 31272 5592 31278
rect 5540 31214 5592 31220
rect 5448 30864 5500 30870
rect 5448 30806 5500 30812
rect 4988 30728 5040 30734
rect 4988 30670 5040 30676
rect 4804 30388 4856 30394
rect 4804 30330 4856 30336
rect 4356 29702 4476 29730
rect 4344 29640 4396 29646
rect 4344 29582 4396 29588
rect 4356 29102 4384 29582
rect 4252 29096 4304 29102
rect 4252 29038 4304 29044
rect 4344 29096 4396 29102
rect 4344 29038 4396 29044
rect 4264 28762 4292 29038
rect 4252 28756 4304 28762
rect 4252 28698 4304 28704
rect 3884 28620 3936 28626
rect 3884 28562 3936 28568
rect 3332 28212 3384 28218
rect 3332 28154 3384 28160
rect 4264 27674 4292 28698
rect 4356 27946 4384 29038
rect 4448 28218 4476 29702
rect 5000 29646 5028 30670
rect 4988 29640 5040 29646
rect 4988 29582 5040 29588
rect 4436 28212 4488 28218
rect 4436 28154 4488 28160
rect 4344 27940 4396 27946
rect 4344 27882 4396 27888
rect 4252 27668 4304 27674
rect 4252 27610 4304 27616
rect 3332 26784 3384 26790
rect 3332 26726 3384 26732
rect 3240 25900 3292 25906
rect 3240 25842 3292 25848
rect 2964 25424 3016 25430
rect 2964 25366 3016 25372
rect 2976 25294 3004 25366
rect 3344 25362 3372 26726
rect 4356 26382 4384 27882
rect 4448 26450 4476 28154
rect 5000 27470 5028 29582
rect 5460 29238 5488 30806
rect 5632 30796 5684 30802
rect 5632 30738 5684 30744
rect 5644 29850 5672 30738
rect 5736 30666 5764 31690
rect 6491 31580 6787 31600
rect 6547 31578 6571 31580
rect 6627 31578 6651 31580
rect 6707 31578 6731 31580
rect 6569 31526 6571 31578
rect 6633 31526 6645 31578
rect 6707 31526 6709 31578
rect 6547 31524 6571 31526
rect 6627 31524 6651 31526
rect 6707 31524 6731 31526
rect 6491 31504 6787 31524
rect 5908 31136 5960 31142
rect 5908 31078 5960 31084
rect 5920 30802 5948 31078
rect 6840 30938 6868 31894
rect 7208 31686 7236 34546
rect 8220 34406 8248 34954
rect 8404 34746 8432 35090
rect 12532 35012 12584 35018
rect 12532 34954 12584 34960
rect 8484 34944 8536 34950
rect 8484 34886 8536 34892
rect 8668 34944 8720 34950
rect 8668 34886 8720 34892
rect 8496 34746 8524 34886
rect 8392 34740 8444 34746
rect 8392 34682 8444 34688
rect 8484 34740 8536 34746
rect 8484 34682 8536 34688
rect 8208 34400 8260 34406
rect 8208 34342 8260 34348
rect 8220 33658 8248 34342
rect 8208 33652 8260 33658
rect 8208 33594 8260 33600
rect 8680 33454 8708 34886
rect 9680 34672 9732 34678
rect 9680 34614 9732 34620
rect 9692 34490 9720 34614
rect 12544 34610 12572 34954
rect 12532 34604 12584 34610
rect 12532 34546 12584 34552
rect 9600 34462 9720 34490
rect 9956 34536 10008 34542
rect 9956 34478 10008 34484
rect 10508 34536 10560 34542
rect 10508 34478 10560 34484
rect 8668 33448 8720 33454
rect 8668 33390 8720 33396
rect 8944 33448 8996 33454
rect 8944 33390 8996 33396
rect 9496 33448 9548 33454
rect 9496 33390 9548 33396
rect 7748 33312 7800 33318
rect 7748 33254 7800 33260
rect 8576 33312 8628 33318
rect 8576 33254 8628 33260
rect 8760 33312 8812 33318
rect 8760 33254 8812 33260
rect 7760 33114 7788 33254
rect 7656 33108 7708 33114
rect 7656 33050 7708 33056
rect 7748 33108 7800 33114
rect 7748 33050 7800 33056
rect 7668 32994 7696 33050
rect 7668 32966 7880 32994
rect 7472 32428 7524 32434
rect 7472 32370 7524 32376
rect 7288 32224 7340 32230
rect 7288 32166 7340 32172
rect 7380 32224 7432 32230
rect 7380 32166 7432 32172
rect 7300 31958 7328 32166
rect 7392 32026 7420 32166
rect 7380 32020 7432 32026
rect 7380 31962 7432 31968
rect 7288 31952 7340 31958
rect 7288 31894 7340 31900
rect 7196 31680 7248 31686
rect 7196 31622 7248 31628
rect 7104 31136 7156 31142
rect 7104 31078 7156 31084
rect 6828 30932 6880 30938
rect 6828 30874 6880 30880
rect 7116 30802 7144 31078
rect 5908 30796 5960 30802
rect 5908 30738 5960 30744
rect 7104 30796 7156 30802
rect 7104 30738 7156 30744
rect 7012 30728 7064 30734
rect 7012 30670 7064 30676
rect 5724 30660 5776 30666
rect 5724 30602 5776 30608
rect 6491 30492 6787 30512
rect 6547 30490 6571 30492
rect 6627 30490 6651 30492
rect 6707 30490 6731 30492
rect 6569 30438 6571 30490
rect 6633 30438 6645 30490
rect 6707 30438 6709 30490
rect 6547 30436 6571 30438
rect 6627 30436 6651 30438
rect 6707 30436 6731 30438
rect 6491 30416 6787 30436
rect 7024 30326 7052 30670
rect 7012 30320 7064 30326
rect 7012 30262 7064 30268
rect 5724 30116 5776 30122
rect 5724 30058 5776 30064
rect 5632 29844 5684 29850
rect 5632 29786 5684 29792
rect 5736 29714 5764 30058
rect 5724 29708 5776 29714
rect 5724 29650 5776 29656
rect 5908 29708 5960 29714
rect 5908 29650 5960 29656
rect 5448 29232 5500 29238
rect 5448 29174 5500 29180
rect 5736 29102 5764 29650
rect 5724 29096 5776 29102
rect 5724 29038 5776 29044
rect 5540 29028 5592 29034
rect 5540 28970 5592 28976
rect 5080 28960 5132 28966
rect 5080 28902 5132 28908
rect 5092 28694 5120 28902
rect 5080 28688 5132 28694
rect 5080 28630 5132 28636
rect 5552 28218 5580 28970
rect 5736 28762 5764 29038
rect 5724 28756 5776 28762
rect 5724 28698 5776 28704
rect 5920 28558 5948 29650
rect 6491 29404 6787 29424
rect 6547 29402 6571 29404
rect 6627 29402 6651 29404
rect 6707 29402 6731 29404
rect 6569 29350 6571 29402
rect 6633 29350 6645 29402
rect 6707 29350 6709 29402
rect 6547 29348 6571 29350
rect 6627 29348 6651 29350
rect 6707 29348 6731 29350
rect 6491 29328 6787 29348
rect 7208 29170 7236 31622
rect 7392 31278 7420 31962
rect 7380 31272 7432 31278
rect 7380 31214 7432 31220
rect 7484 30258 7512 32370
rect 7472 30252 7524 30258
rect 7472 30194 7524 30200
rect 7196 29164 7248 29170
rect 7196 29106 7248 29112
rect 6828 29028 6880 29034
rect 6828 28970 6880 28976
rect 5908 28552 5960 28558
rect 5908 28494 5960 28500
rect 5540 28212 5592 28218
rect 5540 28154 5592 28160
rect 4988 27464 5040 27470
rect 4988 27406 5040 27412
rect 4528 27328 4580 27334
rect 4528 27270 4580 27276
rect 4540 26926 4568 27270
rect 4528 26920 4580 26926
rect 4528 26862 4580 26868
rect 5000 26858 5028 27406
rect 4896 26852 4948 26858
rect 4896 26794 4948 26800
rect 4988 26852 5040 26858
rect 4988 26794 5040 26800
rect 4908 26586 4936 26794
rect 4896 26580 4948 26586
rect 4896 26522 4948 26528
rect 4436 26444 4488 26450
rect 4436 26386 4488 26392
rect 4344 26376 4396 26382
rect 4344 26318 4396 26324
rect 3332 25356 3384 25362
rect 3332 25298 3384 25304
rect 2780 25288 2832 25294
rect 2964 25288 3016 25294
rect 2780 25230 2832 25236
rect 2884 25236 2964 25242
rect 2884 25230 3016 25236
rect 2884 25214 3004 25230
rect 2136 24608 2188 24614
rect 2136 24550 2188 24556
rect 2148 24274 2176 24550
rect 2884 24342 2912 25214
rect 2964 25152 3016 25158
rect 2964 25094 3016 25100
rect 2976 24682 3004 25094
rect 2964 24676 3016 24682
rect 2964 24618 3016 24624
rect 3332 24608 3384 24614
rect 3332 24550 3384 24556
rect 2872 24336 2924 24342
rect 2872 24278 2924 24284
rect 2136 24268 2188 24274
rect 2136 24210 2188 24216
rect 2884 24154 2912 24278
rect 3344 24274 3372 24550
rect 4356 24274 4384 26318
rect 5000 25702 5028 26794
rect 5920 26790 5948 28494
rect 6276 28416 6328 28422
rect 6276 28358 6328 28364
rect 6288 28014 6316 28358
rect 6491 28316 6787 28336
rect 6547 28314 6571 28316
rect 6627 28314 6651 28316
rect 6707 28314 6731 28316
rect 6569 28262 6571 28314
rect 6633 28262 6645 28314
rect 6707 28262 6709 28314
rect 6547 28260 6571 28262
rect 6627 28260 6651 28262
rect 6707 28260 6731 28262
rect 6491 28240 6787 28260
rect 6276 28008 6328 28014
rect 6276 27950 6328 27956
rect 6092 27396 6144 27402
rect 6092 27338 6144 27344
rect 6104 26994 6132 27338
rect 6491 27228 6787 27248
rect 6547 27226 6571 27228
rect 6627 27226 6651 27228
rect 6707 27226 6731 27228
rect 6569 27174 6571 27226
rect 6633 27174 6645 27226
rect 6707 27174 6709 27226
rect 6547 27172 6571 27174
rect 6627 27172 6651 27174
rect 6707 27172 6731 27174
rect 6491 27152 6787 27172
rect 6092 26988 6144 26994
rect 6092 26930 6144 26936
rect 5908 26784 5960 26790
rect 5908 26726 5960 26732
rect 5920 26450 5948 26726
rect 5080 26444 5132 26450
rect 5080 26386 5132 26392
rect 5908 26444 5960 26450
rect 5908 26386 5960 26392
rect 5092 25838 5120 26386
rect 5540 26376 5592 26382
rect 5540 26318 5592 26324
rect 5552 26042 5580 26318
rect 6491 26140 6787 26160
rect 6547 26138 6571 26140
rect 6627 26138 6651 26140
rect 6707 26138 6731 26140
rect 6569 26086 6571 26138
rect 6633 26086 6645 26138
rect 6707 26086 6709 26138
rect 6547 26084 6571 26086
rect 6627 26084 6651 26086
rect 6707 26084 6731 26086
rect 6491 26064 6787 26084
rect 5540 26036 5592 26042
rect 5540 25978 5592 25984
rect 5080 25832 5132 25838
rect 5080 25774 5132 25780
rect 5264 25832 5316 25838
rect 5264 25774 5316 25780
rect 4988 25696 5040 25702
rect 4988 25638 5040 25644
rect 4896 25356 4948 25362
rect 4896 25298 4948 25304
rect 4436 25152 4488 25158
rect 4436 25094 4488 25100
rect 4448 24750 4476 25094
rect 4908 24954 4936 25298
rect 4896 24948 4948 24954
rect 4896 24890 4948 24896
rect 4436 24744 4488 24750
rect 4436 24686 4488 24692
rect 5000 24698 5028 25638
rect 5092 24818 5120 25774
rect 5276 25498 5304 25774
rect 5264 25492 5316 25498
rect 5264 25434 5316 25440
rect 5172 25288 5224 25294
rect 5172 25230 5224 25236
rect 5080 24812 5132 24818
rect 5080 24754 5132 24760
rect 5000 24682 5120 24698
rect 5000 24676 5132 24682
rect 5000 24670 5080 24676
rect 5080 24618 5132 24624
rect 5092 24426 5120 24618
rect 5184 24614 5212 25230
rect 5172 24608 5224 24614
rect 5172 24550 5224 24556
rect 5092 24398 5212 24426
rect 5184 24274 5212 24398
rect 3332 24268 3384 24274
rect 3332 24210 3384 24216
rect 4344 24268 4396 24274
rect 4344 24210 4396 24216
rect 5172 24268 5224 24274
rect 5172 24210 5224 24216
rect 2884 24126 3004 24154
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 2780 24064 2832 24070
rect 2832 24012 2912 24018
rect 2780 24006 2912 24012
rect 2792 23990 2912 24006
rect 2688 23248 2740 23254
rect 2688 23190 2740 23196
rect 2700 22710 2728 23190
rect 2688 22704 2740 22710
rect 2608 22652 2688 22658
rect 2608 22646 2740 22652
rect 2608 22630 2728 22646
rect 1676 21888 1728 21894
rect 1676 21830 1728 21836
rect 1688 21554 1716 21830
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 2608 21350 2636 22630
rect 2688 22568 2740 22574
rect 2688 22510 2740 22516
rect 2700 22166 2728 22510
rect 2780 22432 2832 22438
rect 2780 22374 2832 22380
rect 2688 22160 2740 22166
rect 2688 22102 2740 22108
rect 2596 21344 2648 21350
rect 2596 21286 2648 21292
rect 1766 20496 1822 20505
rect 1766 20431 1768 20440
rect 1820 20431 1822 20440
rect 1768 20402 1820 20408
rect 1952 20324 2004 20330
rect 1952 20266 2004 20272
rect 1964 19786 1992 20266
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 1952 19780 2004 19786
rect 1952 19722 2004 19728
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1688 19378 1716 19654
rect 1676 19372 1728 19378
rect 1676 19314 1728 19320
rect 2240 18970 2268 19790
rect 2608 19258 2636 21286
rect 2700 19922 2728 22102
rect 2792 22030 2820 22374
rect 2780 22024 2832 22030
rect 2780 21966 2832 21972
rect 2688 19916 2740 19922
rect 2688 19858 2740 19864
rect 2424 19242 2636 19258
rect 2412 19236 2636 19242
rect 2464 19230 2636 19236
rect 2412 19178 2464 19184
rect 2228 18964 2280 18970
rect 2228 18906 2280 18912
rect 2700 18902 2728 19858
rect 2688 18896 2740 18902
rect 2688 18838 2740 18844
rect 2504 18216 2556 18222
rect 2504 18158 2556 18164
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 2516 17882 2544 18158
rect 2504 17876 2556 17882
rect 2504 17818 2556 17824
rect 2596 17740 2648 17746
rect 2596 17682 2648 17688
rect 2608 17542 2636 17682
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2608 17134 2636 17478
rect 2792 17338 2820 18158
rect 2884 17882 2912 23990
rect 2976 23866 3004 24126
rect 3792 24132 3844 24138
rect 3792 24074 3844 24080
rect 2964 23860 3016 23866
rect 2964 23802 3016 23808
rect 3332 23588 3384 23594
rect 3332 23530 3384 23536
rect 2964 23180 3016 23186
rect 2964 23122 3016 23128
rect 2976 22574 3004 23122
rect 3344 22778 3372 23530
rect 3332 22772 3384 22778
rect 3332 22714 3384 22720
rect 2964 22568 3016 22574
rect 2964 22510 3016 22516
rect 3332 22568 3384 22574
rect 3332 22510 3384 22516
rect 2976 22094 3004 22510
rect 3344 22166 3372 22510
rect 3332 22160 3384 22166
rect 3332 22102 3384 22108
rect 2976 22066 3096 22094
rect 2964 21888 3016 21894
rect 2964 21830 3016 21836
rect 2976 20874 3004 21830
rect 3068 21486 3096 22066
rect 3056 21480 3108 21486
rect 3056 21422 3108 21428
rect 3148 21004 3200 21010
rect 3148 20946 3200 20952
rect 3332 21004 3384 21010
rect 3332 20946 3384 20952
rect 2964 20868 3016 20874
rect 2964 20810 3016 20816
rect 3160 20602 3188 20946
rect 3344 20602 3372 20946
rect 3148 20596 3200 20602
rect 3148 20538 3200 20544
rect 3332 20596 3384 20602
rect 3332 20538 3384 20544
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 3068 18154 3096 19994
rect 3160 19718 3188 20538
rect 3344 20058 3372 20538
rect 3332 20052 3384 20058
rect 3332 19994 3384 20000
rect 3332 19916 3384 19922
rect 3332 19858 3384 19864
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3344 19514 3372 19858
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 3344 18834 3372 19450
rect 3332 18828 3384 18834
rect 3332 18770 3384 18776
rect 3240 18216 3292 18222
rect 3240 18158 3292 18164
rect 3056 18148 3108 18154
rect 3056 18090 3108 18096
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 3068 17814 3096 18090
rect 3056 17808 3108 17814
rect 3056 17750 3108 17756
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2596 17128 2648 17134
rect 2596 17070 2648 17076
rect 2884 17066 2912 17614
rect 2872 17060 2924 17066
rect 2872 17002 2924 17008
rect 1676 15972 1728 15978
rect 1676 15914 1728 15920
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 1688 15706 1716 15914
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 2700 15638 2728 15914
rect 2688 15632 2740 15638
rect 2688 15574 2740 15580
rect 2700 14890 2728 15574
rect 2884 15314 2912 17002
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 2976 15502 3004 16594
rect 3056 16448 3108 16454
rect 3056 16390 3108 16396
rect 3068 15570 3096 16390
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2884 15286 3004 15314
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1780 12850 1808 13126
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 1768 12368 1820 12374
rect 1766 12336 1768 12345
rect 1820 12336 1822 12345
rect 1766 12271 1822 12280
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1780 11218 1808 11494
rect 2700 11286 2728 12582
rect 2884 12442 2912 13330
rect 2976 13326 3004 15286
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 2976 12986 3004 13262
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2976 11830 3004 12174
rect 2964 11824 3016 11830
rect 2964 11766 3016 11772
rect 2688 11280 2740 11286
rect 2688 11222 2740 11228
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2792 10266 2820 10950
rect 2884 10674 2912 11086
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1780 9586 1808 9862
rect 2884 9722 2912 9998
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 2320 9444 2372 9450
rect 2320 9386 2372 9392
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 2332 8022 2360 9386
rect 2884 9042 2912 9658
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2976 8974 3004 11766
rect 3068 11694 3096 13262
rect 3252 12238 3280 18158
rect 3424 16720 3476 16726
rect 3424 16662 3476 16668
rect 3332 16652 3384 16658
rect 3332 16594 3384 16600
rect 3344 15042 3372 16594
rect 3436 16114 3464 16662
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 3436 15570 3464 16050
rect 3424 15564 3476 15570
rect 3424 15506 3476 15512
rect 3436 15094 3464 15125
rect 3424 15088 3476 15094
rect 3344 15036 3424 15042
rect 3344 15030 3476 15036
rect 3344 15014 3464 15030
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 3344 14346 3372 14894
rect 3436 14618 3464 15014
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3332 14340 3384 14346
rect 3332 14282 3384 14288
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3068 11150 3096 11630
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 3068 10810 3096 11086
rect 3436 11014 3464 11630
rect 3424 11008 3476 11014
rect 3424 10950 3476 10956
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3344 10062 3372 10542
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3344 9450 3372 9998
rect 3804 9518 3832 24074
rect 4356 23798 4384 24210
rect 4528 24200 4580 24206
rect 4528 24142 4580 24148
rect 4344 23792 4396 23798
rect 4344 23734 4396 23740
rect 4436 23724 4488 23730
rect 4436 23666 4488 23672
rect 4160 23112 4212 23118
rect 4160 23054 4212 23060
rect 4172 22778 4200 23054
rect 4160 22772 4212 22778
rect 4160 22714 4212 22720
rect 4448 22574 4476 23666
rect 4344 22568 4396 22574
rect 4344 22510 4396 22516
rect 4436 22568 4488 22574
rect 4436 22510 4488 22516
rect 4252 22160 4304 22166
rect 4252 22102 4304 22108
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 4080 21486 4108 21966
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 3884 21480 3936 21486
rect 3884 21422 3936 21428
rect 4068 21480 4120 21486
rect 4068 21422 4120 21428
rect 3896 20890 3924 21422
rect 3976 21344 4028 21350
rect 3976 21286 4028 21292
rect 3988 21078 4016 21286
rect 3976 21072 4028 21078
rect 3976 21014 4028 21020
rect 3896 20862 4016 20890
rect 3988 20806 4016 20862
rect 3976 20800 4028 20806
rect 3976 20742 4028 20748
rect 3988 20466 4016 20742
rect 4080 20602 4108 21422
rect 4068 20596 4120 20602
rect 4068 20538 4120 20544
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 3884 20392 3936 20398
rect 3884 20334 3936 20340
rect 3896 19922 3924 20334
rect 3884 19916 3936 19922
rect 3884 19858 3936 19864
rect 3988 19514 4016 20402
rect 4080 19718 4108 20538
rect 4172 20058 4200 21490
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 4172 19174 4200 19994
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 4172 18902 4200 19110
rect 4160 18896 4212 18902
rect 4160 18838 4212 18844
rect 4068 18692 4120 18698
rect 4068 18634 4120 18640
rect 3884 18080 3936 18086
rect 3884 18022 3936 18028
rect 3896 12374 3924 18022
rect 4080 16425 4108 18634
rect 4264 18154 4292 22102
rect 4356 21146 4384 22510
rect 4540 21332 4568 24142
rect 4620 24132 4672 24138
rect 4620 24074 4672 24080
rect 4632 23730 4660 24074
rect 4620 23724 4672 23730
rect 4620 23666 4672 23672
rect 4632 22098 4660 23666
rect 4896 23656 4948 23662
rect 4896 23598 4948 23604
rect 4908 23050 4936 23598
rect 5184 23254 5212 24210
rect 5276 23662 5304 25434
rect 5552 25430 5580 25978
rect 5540 25424 5592 25430
rect 5540 25366 5592 25372
rect 5632 25152 5684 25158
rect 5632 25094 5684 25100
rect 5644 24818 5672 25094
rect 6491 25052 6787 25072
rect 6547 25050 6571 25052
rect 6627 25050 6651 25052
rect 6707 25050 6731 25052
rect 6569 24998 6571 25050
rect 6633 24998 6645 25050
rect 6707 24998 6709 25050
rect 6547 24996 6571 24998
rect 6627 24996 6651 24998
rect 6707 24996 6731 24998
rect 6491 24976 6787 24996
rect 5632 24812 5684 24818
rect 5632 24754 5684 24760
rect 6276 24336 6328 24342
rect 6276 24278 6328 24284
rect 5264 23656 5316 23662
rect 5264 23598 5316 23604
rect 5172 23248 5224 23254
rect 5172 23190 5224 23196
rect 4896 23044 4948 23050
rect 4896 22986 4948 22992
rect 4712 22976 4764 22982
rect 4712 22918 4764 22924
rect 4724 22658 4752 22918
rect 4724 22642 4844 22658
rect 4712 22636 4844 22642
rect 4764 22630 4844 22636
rect 4712 22578 4764 22584
rect 4712 22500 4764 22506
rect 4712 22442 4764 22448
rect 4724 22234 4752 22442
rect 4712 22228 4764 22234
rect 4712 22170 4764 22176
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 4816 21554 4844 22630
rect 4908 22098 4936 22986
rect 4896 22092 4948 22098
rect 4896 22034 4948 22040
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 5000 21554 5028 21830
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 4988 21548 5040 21554
rect 4988 21490 5040 21496
rect 4540 21304 4660 21332
rect 4344 21140 4396 21146
rect 4344 21082 4396 21088
rect 4436 20936 4488 20942
rect 4436 20878 4488 20884
rect 4528 20936 4580 20942
rect 4528 20878 4580 20884
rect 4448 19514 4476 20878
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 4540 19310 4568 20878
rect 4632 20874 4660 21304
rect 4620 20868 4672 20874
rect 4620 20810 4672 20816
rect 4816 20398 4844 21490
rect 4804 20392 4856 20398
rect 4724 20352 4804 20380
rect 4724 19854 4752 20352
rect 4804 20334 4856 20340
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 5092 19922 5120 20198
rect 5276 19990 5304 23598
rect 5356 23112 5408 23118
rect 5356 23054 5408 23060
rect 5816 23112 5868 23118
rect 5816 23054 5868 23060
rect 5368 22098 5396 23054
rect 5828 22710 5856 23054
rect 5816 22704 5868 22710
rect 5816 22646 5868 22652
rect 6288 22574 6316 24278
rect 6491 23964 6787 23984
rect 6547 23962 6571 23964
rect 6627 23962 6651 23964
rect 6707 23962 6731 23964
rect 6569 23910 6571 23962
rect 6633 23910 6645 23962
rect 6707 23910 6709 23962
rect 6547 23908 6571 23910
rect 6627 23908 6651 23910
rect 6707 23908 6731 23910
rect 6491 23888 6787 23908
rect 6491 22876 6787 22896
rect 6547 22874 6571 22876
rect 6627 22874 6651 22876
rect 6707 22874 6731 22876
rect 6569 22822 6571 22874
rect 6633 22822 6645 22874
rect 6707 22822 6709 22874
rect 6547 22820 6571 22822
rect 6627 22820 6651 22822
rect 6707 22820 6731 22822
rect 6491 22800 6787 22820
rect 6276 22568 6328 22574
rect 6276 22510 6328 22516
rect 6736 22432 6788 22438
rect 6736 22374 6788 22380
rect 6748 22166 6776 22374
rect 6736 22160 6788 22166
rect 6736 22102 6788 22108
rect 5356 22092 5408 22098
rect 5356 22034 5408 22040
rect 5540 22092 5592 22098
rect 5540 22034 5592 22040
rect 5552 21010 5580 22034
rect 6491 21788 6787 21808
rect 6547 21786 6571 21788
rect 6627 21786 6651 21788
rect 6707 21786 6731 21788
rect 6569 21734 6571 21786
rect 6633 21734 6645 21786
rect 6707 21734 6709 21786
rect 6547 21732 6571 21734
rect 6627 21732 6651 21734
rect 6707 21732 6731 21734
rect 6491 21712 6787 21732
rect 5724 21344 5776 21350
rect 5724 21286 5776 21292
rect 5448 21004 5500 21010
rect 5448 20946 5500 20952
rect 5540 21004 5592 21010
rect 5540 20946 5592 20952
rect 5460 20398 5488 20946
rect 5736 20398 5764 21286
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 6380 20806 6408 20946
rect 6368 20800 6420 20806
rect 6368 20742 6420 20748
rect 5448 20392 5500 20398
rect 5448 20334 5500 20340
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 5460 20058 5488 20334
rect 5448 20052 5500 20058
rect 5448 19994 5500 20000
rect 5264 19984 5316 19990
rect 5264 19926 5316 19932
rect 5080 19916 5132 19922
rect 5080 19858 5132 19864
rect 5632 19916 5684 19922
rect 5632 19858 5684 19864
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 4724 19310 4752 19790
rect 5092 19310 5120 19858
rect 5644 19378 5672 19858
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 4528 19304 4580 19310
rect 4528 19246 4580 19252
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 4540 18970 4568 19246
rect 4528 18964 4580 18970
rect 4528 18906 4580 18912
rect 5092 18902 5120 19246
rect 5552 18970 5580 19246
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5080 18896 5132 18902
rect 5080 18838 5132 18844
rect 5092 18290 5120 18838
rect 5724 18828 5776 18834
rect 5724 18770 5776 18776
rect 6184 18828 6236 18834
rect 6184 18770 6236 18776
rect 5736 18630 5764 18770
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5080 18284 5132 18290
rect 5080 18226 5132 18232
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 4252 18148 4304 18154
rect 4252 18090 4304 18096
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4172 16658 4200 18022
rect 4264 17134 4292 18090
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 4712 17808 4764 17814
rect 4712 17750 4764 17756
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4252 17128 4304 17134
rect 4252 17070 4304 17076
rect 4356 16794 4384 17682
rect 4724 17338 4752 17750
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 4908 17338 4936 17478
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 4896 17332 4948 17338
rect 4896 17274 4948 17280
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 4344 16788 4396 16794
rect 4344 16730 4396 16736
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 4066 16416 4122 16425
rect 4066 16351 4122 16360
rect 4172 16130 4200 16594
rect 4816 16250 4844 17070
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4172 16102 4292 16130
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 4080 15026 4108 15438
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4080 14618 4108 14962
rect 4172 14890 4200 15982
rect 4264 14958 4292 16102
rect 4528 15360 4580 15366
rect 4528 15302 4580 15308
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 4540 14890 4568 15302
rect 4160 14884 4212 14890
rect 4160 14826 4212 14832
rect 4528 14884 4580 14890
rect 4528 14826 4580 14832
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4172 14550 4200 14826
rect 4540 14550 4568 14826
rect 4160 14544 4212 14550
rect 4160 14486 4212 14492
rect 4528 14544 4580 14550
rect 4528 14486 4580 14492
rect 4172 14346 4200 14486
rect 4160 14340 4212 14346
rect 4160 14282 4212 14288
rect 5000 13734 5028 18022
rect 5276 17814 5304 18158
rect 6196 18154 6224 18770
rect 6184 18148 6236 18154
rect 6184 18090 6236 18096
rect 5264 17808 5316 17814
rect 5264 17750 5316 17756
rect 6196 17746 6224 18090
rect 6380 17746 6408 20742
rect 6491 20700 6787 20720
rect 6547 20698 6571 20700
rect 6627 20698 6651 20700
rect 6707 20698 6731 20700
rect 6569 20646 6571 20698
rect 6633 20646 6645 20698
rect 6707 20646 6709 20698
rect 6547 20644 6571 20646
rect 6627 20644 6651 20646
rect 6707 20644 6731 20646
rect 6491 20624 6787 20644
rect 6840 20058 6868 28970
rect 7208 26382 7236 29106
rect 7484 28558 7512 30194
rect 7656 29640 7708 29646
rect 7656 29582 7708 29588
rect 7668 29238 7696 29582
rect 7656 29232 7708 29238
rect 7656 29174 7708 29180
rect 7668 29102 7696 29174
rect 7656 29096 7708 29102
rect 7656 29038 7708 29044
rect 7472 28552 7524 28558
rect 7472 28494 7524 28500
rect 7288 27328 7340 27334
rect 7340 27288 7420 27316
rect 7288 27270 7340 27276
rect 7196 26376 7248 26382
rect 7196 26318 7248 26324
rect 7208 25974 7236 26318
rect 7196 25968 7248 25974
rect 7196 25910 7248 25916
rect 7012 25424 7064 25430
rect 7012 25366 7064 25372
rect 6920 24268 6972 24274
rect 6920 24210 6972 24216
rect 6932 23662 6960 24210
rect 6920 23656 6972 23662
rect 6920 23598 6972 23604
rect 6932 22778 6960 23598
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6932 22098 6960 22714
rect 7024 22642 7052 25366
rect 7104 25288 7156 25294
rect 7104 25230 7156 25236
rect 7116 24954 7144 25230
rect 7104 24948 7156 24954
rect 7104 24890 7156 24896
rect 7208 24750 7236 25910
rect 7288 25900 7340 25906
rect 7288 25842 7340 25848
rect 7300 24954 7328 25842
rect 7392 25770 7420 27288
rect 7472 26784 7524 26790
rect 7472 26726 7524 26732
rect 7484 26586 7512 26726
rect 7472 26580 7524 26586
rect 7472 26522 7524 26528
rect 7484 25906 7512 26522
rect 7852 26330 7880 32966
rect 8300 32972 8352 32978
rect 8300 32914 8352 32920
rect 8312 32570 8340 32914
rect 8484 32768 8536 32774
rect 8484 32710 8536 32716
rect 8300 32564 8352 32570
rect 8300 32506 8352 32512
rect 8496 32366 8524 32710
rect 8588 32570 8616 33254
rect 8576 32564 8628 32570
rect 8576 32506 8628 32512
rect 8484 32360 8536 32366
rect 8484 32302 8536 32308
rect 8772 32298 8800 33254
rect 8956 32774 8984 33390
rect 8944 32768 8996 32774
rect 8944 32710 8996 32716
rect 8760 32292 8812 32298
rect 8760 32234 8812 32240
rect 8208 31136 8260 31142
rect 8208 31078 8260 31084
rect 8220 30190 8248 31078
rect 8208 30184 8260 30190
rect 8208 30126 8260 30132
rect 8024 29708 8076 29714
rect 8024 29650 8076 29656
rect 8036 29306 8064 29650
rect 8024 29300 8076 29306
rect 8024 29242 8076 29248
rect 8220 29170 8248 30126
rect 8576 30048 8628 30054
rect 8576 29990 8628 29996
rect 8588 29714 8616 29990
rect 8576 29708 8628 29714
rect 8576 29650 8628 29656
rect 8208 29164 8260 29170
rect 8208 29106 8260 29112
rect 8588 28626 8616 29650
rect 8852 28960 8904 28966
rect 8852 28902 8904 28908
rect 8864 28762 8892 28902
rect 8852 28756 8904 28762
rect 8852 28698 8904 28704
rect 8300 28620 8352 28626
rect 8300 28562 8352 28568
rect 8576 28620 8628 28626
rect 8576 28562 8628 28568
rect 8208 28008 8260 28014
rect 8312 27996 8340 28562
rect 8260 27968 8340 27996
rect 8208 27950 8260 27956
rect 8208 27872 8260 27878
rect 8208 27814 8260 27820
rect 7932 26988 7984 26994
rect 7932 26930 7984 26936
rect 7944 26450 7972 26930
rect 8220 26926 8248 27814
rect 8208 26920 8260 26926
rect 8208 26862 8260 26868
rect 7932 26444 7984 26450
rect 7932 26386 7984 26392
rect 7852 26302 7972 26330
rect 7840 26240 7892 26246
rect 7840 26182 7892 26188
rect 7472 25900 7524 25906
rect 7472 25842 7524 25848
rect 7852 25838 7880 26182
rect 7840 25832 7892 25838
rect 7840 25774 7892 25780
rect 7380 25764 7432 25770
rect 7380 25706 7432 25712
rect 7392 25362 7420 25706
rect 7472 25696 7524 25702
rect 7472 25638 7524 25644
rect 7380 25356 7432 25362
rect 7380 25298 7432 25304
rect 7484 25226 7512 25638
rect 7944 25362 7972 26302
rect 8312 25498 8340 27968
rect 8392 28008 8444 28014
rect 8392 27950 8444 27956
rect 8404 27538 8432 27950
rect 8392 27532 8444 27538
rect 8392 27474 8444 27480
rect 8404 26586 8432 27474
rect 8760 27464 8812 27470
rect 8760 27406 8812 27412
rect 8668 26920 8720 26926
rect 8668 26862 8720 26868
rect 8392 26580 8444 26586
rect 8392 26522 8444 26528
rect 8680 26042 8708 26862
rect 8772 26790 8800 27406
rect 8956 26926 8984 32710
rect 9128 29504 9180 29510
rect 9128 29446 9180 29452
rect 9140 28762 9168 29446
rect 9508 29102 9536 33390
rect 9600 32774 9628 34462
rect 9680 33992 9732 33998
rect 9680 33934 9732 33940
rect 9692 32910 9720 33934
rect 9968 33386 9996 34478
rect 10140 34400 10192 34406
rect 10140 34342 10192 34348
rect 10152 34134 10180 34342
rect 10140 34128 10192 34134
rect 10140 34070 10192 34076
rect 10416 33448 10468 33454
rect 10416 33390 10468 33396
rect 9956 33380 10008 33386
rect 9956 33322 10008 33328
rect 9968 32910 9996 33322
rect 10428 32978 10456 33390
rect 10520 33114 10548 34478
rect 12440 34400 12492 34406
rect 12440 34342 12492 34348
rect 12532 34400 12584 34406
rect 12532 34342 12584 34348
rect 12026 34300 12322 34320
rect 12082 34298 12106 34300
rect 12162 34298 12186 34300
rect 12242 34298 12266 34300
rect 12104 34246 12106 34298
rect 12168 34246 12180 34298
rect 12242 34246 12244 34298
rect 12082 34244 12106 34246
rect 12162 34244 12186 34246
rect 12242 34244 12266 34246
rect 12026 34224 12322 34244
rect 12452 34202 12480 34342
rect 12544 34202 12572 34342
rect 12440 34196 12492 34202
rect 12440 34138 12492 34144
rect 12532 34196 12584 34202
rect 12532 34138 12584 34144
rect 11244 33856 11296 33862
rect 11244 33798 11296 33804
rect 11256 33318 11284 33798
rect 12544 33658 12572 34138
rect 12532 33652 12584 33658
rect 12532 33594 12584 33600
rect 12532 33448 12584 33454
rect 12532 33390 12584 33396
rect 11244 33312 11296 33318
rect 11244 33254 11296 33260
rect 10508 33108 10560 33114
rect 10508 33050 10560 33056
rect 11256 32978 11284 33254
rect 12026 33212 12322 33232
rect 12082 33210 12106 33212
rect 12162 33210 12186 33212
rect 12242 33210 12266 33212
rect 12104 33158 12106 33210
rect 12168 33158 12180 33210
rect 12242 33158 12244 33210
rect 12082 33156 12106 33158
rect 12162 33156 12186 33158
rect 12242 33156 12266 33158
rect 12026 33136 12322 33156
rect 10232 32972 10284 32978
rect 10232 32914 10284 32920
rect 10416 32972 10468 32978
rect 10416 32914 10468 32920
rect 11244 32972 11296 32978
rect 11244 32914 11296 32920
rect 9680 32904 9732 32910
rect 9680 32846 9732 32852
rect 9956 32904 10008 32910
rect 9956 32846 10008 32852
rect 9588 32768 9640 32774
rect 9588 32710 9640 32716
rect 9692 32366 9720 32846
rect 9588 32360 9640 32366
rect 9588 32302 9640 32308
rect 9680 32360 9732 32366
rect 9680 32302 9732 32308
rect 9600 32230 9628 32302
rect 9588 32224 9640 32230
rect 9588 32166 9640 32172
rect 9600 32026 9628 32166
rect 9588 32020 9640 32026
rect 9588 31962 9640 31968
rect 9692 31754 9720 32302
rect 9968 32298 9996 32846
rect 10048 32768 10100 32774
rect 10048 32710 10100 32716
rect 10060 32366 10088 32710
rect 10048 32360 10100 32366
rect 10048 32302 10100 32308
rect 9956 32292 10008 32298
rect 9956 32234 10008 32240
rect 9864 31816 9916 31822
rect 9864 31758 9916 31764
rect 9680 31748 9732 31754
rect 9680 31690 9732 31696
rect 9876 31498 9904 31758
rect 9692 31470 9904 31498
rect 9496 29096 9548 29102
rect 9496 29038 9548 29044
rect 9128 28756 9180 28762
rect 9128 28698 9180 28704
rect 9508 28082 9536 29038
rect 9692 28626 9720 31470
rect 9968 31362 9996 32234
rect 10244 32026 10272 32914
rect 10324 32904 10376 32910
rect 10324 32846 10376 32852
rect 10232 32020 10284 32026
rect 10232 31962 10284 31968
rect 10048 31748 10100 31754
rect 10048 31690 10100 31696
rect 9876 31334 9996 31362
rect 9876 31210 9904 31334
rect 9956 31272 10008 31278
rect 10060 31226 10088 31690
rect 10008 31220 10088 31226
rect 9956 31214 10088 31220
rect 9772 31204 9824 31210
rect 9772 31146 9824 31152
rect 9864 31204 9916 31210
rect 9864 31146 9916 31152
rect 9968 31198 10088 31214
rect 9784 29850 9812 31146
rect 9876 30546 9904 31146
rect 9968 30734 9996 31198
rect 10140 31136 10192 31142
rect 10140 31078 10192 31084
rect 10048 30796 10100 30802
rect 10048 30738 10100 30744
rect 9956 30728 10008 30734
rect 9956 30670 10008 30676
rect 9876 30518 9996 30546
rect 9772 29844 9824 29850
rect 9772 29786 9824 29792
rect 9864 29572 9916 29578
rect 9864 29514 9916 29520
rect 9876 29306 9904 29514
rect 9864 29300 9916 29306
rect 9864 29242 9916 29248
rect 9968 29102 9996 30518
rect 10060 30394 10088 30738
rect 10048 30388 10100 30394
rect 10048 30330 10100 30336
rect 10152 30190 10180 31078
rect 10140 30184 10192 30190
rect 10140 30126 10192 30132
rect 10232 29708 10284 29714
rect 10232 29650 10284 29656
rect 9956 29096 10008 29102
rect 9956 29038 10008 29044
rect 9680 28620 9732 28626
rect 9680 28562 9732 28568
rect 9864 28620 9916 28626
rect 9864 28562 9916 28568
rect 9496 28076 9548 28082
rect 9496 28018 9548 28024
rect 9036 26988 9088 26994
rect 9036 26930 9088 26936
rect 8944 26920 8996 26926
rect 8944 26862 8996 26868
rect 8760 26784 8812 26790
rect 8760 26726 8812 26732
rect 8668 26036 8720 26042
rect 8668 25978 8720 25984
rect 8760 25832 8812 25838
rect 8760 25774 8812 25780
rect 8300 25492 8352 25498
rect 8300 25434 8352 25440
rect 7932 25356 7984 25362
rect 7932 25298 7984 25304
rect 7472 25220 7524 25226
rect 7472 25162 7524 25168
rect 7288 24948 7340 24954
rect 7288 24890 7340 24896
rect 7196 24744 7248 24750
rect 7196 24686 7248 24692
rect 7564 24404 7616 24410
rect 7564 24346 7616 24352
rect 7576 24274 7604 24346
rect 7944 24342 7972 25298
rect 8300 24744 8352 24750
rect 8300 24686 8352 24692
rect 7932 24336 7984 24342
rect 7932 24278 7984 24284
rect 7564 24268 7616 24274
rect 7564 24210 7616 24216
rect 8312 23610 8340 24686
rect 8668 24132 8720 24138
rect 8668 24074 8720 24080
rect 8312 23582 8524 23610
rect 7104 23180 7156 23186
rect 7104 23122 7156 23128
rect 7012 22636 7064 22642
rect 7012 22578 7064 22584
rect 6920 22092 6972 22098
rect 6920 22034 6972 22040
rect 6920 21140 6972 21146
rect 6920 21082 6972 21088
rect 6932 20602 6960 21082
rect 7024 21010 7052 22578
rect 7116 22030 7144 23122
rect 8312 23050 8340 23582
rect 8496 23526 8524 23582
rect 8392 23520 8444 23526
rect 8392 23462 8444 23468
rect 8484 23520 8536 23526
rect 8484 23462 8536 23468
rect 8024 23044 8076 23050
rect 8024 22986 8076 22992
rect 8300 23044 8352 23050
rect 8300 22986 8352 22992
rect 7932 22636 7984 22642
rect 7932 22578 7984 22584
rect 7944 22098 7972 22578
rect 8036 22438 8064 22986
rect 8404 22642 8432 23462
rect 8392 22636 8444 22642
rect 8392 22578 8444 22584
rect 8024 22432 8076 22438
rect 8024 22374 8076 22380
rect 7472 22092 7524 22098
rect 7472 22034 7524 22040
rect 7932 22092 7984 22098
rect 7932 22034 7984 22040
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 7288 21956 7340 21962
rect 7288 21898 7340 21904
rect 7300 21146 7328 21898
rect 7288 21140 7340 21146
rect 7288 21082 7340 21088
rect 7012 21004 7064 21010
rect 7012 20946 7064 20952
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 7024 20330 7052 20946
rect 7012 20324 7064 20330
rect 7012 20266 7064 20272
rect 6828 20052 6880 20058
rect 6828 19994 6880 20000
rect 6491 19612 6787 19632
rect 6547 19610 6571 19612
rect 6627 19610 6651 19612
rect 6707 19610 6731 19612
rect 6569 19558 6571 19610
rect 6633 19558 6645 19610
rect 6707 19558 6709 19610
rect 6547 19556 6571 19558
rect 6627 19556 6651 19558
rect 6707 19556 6731 19558
rect 6491 19536 6787 19556
rect 6840 18834 6868 19994
rect 7024 19242 7052 20266
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 7116 19378 7144 19790
rect 7104 19372 7156 19378
rect 7104 19314 7156 19320
rect 7012 19236 7064 19242
rect 7012 19178 7064 19184
rect 6828 18828 6880 18834
rect 6828 18770 6880 18776
rect 6491 18524 6787 18544
rect 6547 18522 6571 18524
rect 6627 18522 6651 18524
rect 6707 18522 6731 18524
rect 6569 18470 6571 18522
rect 6633 18470 6645 18522
rect 6707 18470 6709 18522
rect 6547 18468 6571 18470
rect 6627 18468 6651 18470
rect 6707 18468 6731 18470
rect 6491 18448 6787 18468
rect 6840 18222 6868 18770
rect 7300 18222 7328 21082
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7484 17746 7512 22034
rect 8036 21486 8064 22374
rect 8680 21486 8708 24074
rect 8772 22642 8800 25774
rect 8852 24608 8904 24614
rect 8852 24550 8904 24556
rect 8864 23866 8892 24550
rect 8852 23860 8904 23866
rect 8852 23802 8904 23808
rect 8760 22636 8812 22642
rect 8760 22578 8812 22584
rect 8772 21486 8800 22578
rect 8024 21480 8076 21486
rect 8024 21422 8076 21428
rect 8668 21480 8720 21486
rect 8668 21422 8720 21428
rect 8760 21480 8812 21486
rect 8760 21422 8812 21428
rect 8208 21344 8260 21350
rect 8208 21286 8260 21292
rect 8220 21078 8248 21286
rect 8680 21146 8708 21422
rect 8668 21140 8720 21146
rect 8668 21082 8720 21088
rect 8208 21072 8260 21078
rect 8208 21014 8260 21020
rect 8208 20936 8260 20942
rect 8208 20878 8260 20884
rect 8220 20602 8248 20878
rect 8392 20800 8444 20806
rect 8392 20742 8444 20748
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 8220 18426 8248 20538
rect 8404 20466 8432 20742
rect 8392 20460 8444 20466
rect 8392 20402 8444 20408
rect 8956 20330 8984 26862
rect 9048 26246 9076 26930
rect 9508 26926 9536 28018
rect 9876 27130 9904 28562
rect 9968 27538 9996 29038
rect 10244 28762 10272 29650
rect 10232 28756 10284 28762
rect 10232 28698 10284 28704
rect 10048 28552 10100 28558
rect 10048 28494 10100 28500
rect 9956 27532 10008 27538
rect 9956 27474 10008 27480
rect 10060 27470 10088 28494
rect 10232 28008 10284 28014
rect 10232 27950 10284 27956
rect 10140 27940 10192 27946
rect 10140 27882 10192 27888
rect 10152 27606 10180 27882
rect 10140 27600 10192 27606
rect 10140 27542 10192 27548
rect 10048 27464 10100 27470
rect 10048 27406 10100 27412
rect 9864 27124 9916 27130
rect 9864 27066 9916 27072
rect 9496 26920 9548 26926
rect 9496 26862 9548 26868
rect 10152 26518 10180 27542
rect 10244 27538 10272 27950
rect 10232 27532 10284 27538
rect 10232 27474 10284 27480
rect 10244 26586 10272 27474
rect 10336 26858 10364 32846
rect 10428 31890 10456 32914
rect 12544 32434 12572 33390
rect 12532 32428 12584 32434
rect 12532 32370 12584 32376
rect 11152 32224 11204 32230
rect 11152 32166 11204 32172
rect 12440 32224 12492 32230
rect 12440 32166 12492 32172
rect 11164 31958 11192 32166
rect 12026 32124 12322 32144
rect 12082 32122 12106 32124
rect 12162 32122 12186 32124
rect 12242 32122 12266 32124
rect 12104 32070 12106 32122
rect 12168 32070 12180 32122
rect 12242 32070 12244 32122
rect 12082 32068 12106 32070
rect 12162 32068 12186 32070
rect 12242 32068 12266 32070
rect 12026 32048 12322 32068
rect 12452 32026 12480 32166
rect 12440 32020 12492 32026
rect 12440 31962 12492 31968
rect 11152 31952 11204 31958
rect 11152 31894 11204 31900
rect 10416 31884 10468 31890
rect 10416 31826 10468 31832
rect 10428 27606 10456 31826
rect 12544 31686 12572 32370
rect 12532 31680 12584 31686
rect 12532 31622 12584 31628
rect 12544 31346 12572 31622
rect 12532 31340 12584 31346
rect 12532 31282 12584 31288
rect 11612 31272 11664 31278
rect 11612 31214 11664 31220
rect 11624 30938 11652 31214
rect 12440 31136 12492 31142
rect 12440 31078 12492 31084
rect 12026 31036 12322 31056
rect 12082 31034 12106 31036
rect 12162 31034 12186 31036
rect 12242 31034 12266 31036
rect 12104 30982 12106 31034
rect 12168 30982 12180 31034
rect 12242 30982 12244 31034
rect 12082 30980 12106 30982
rect 12162 30980 12186 30982
rect 12242 30980 12266 30982
rect 12026 30960 12322 30980
rect 12452 30938 12480 31078
rect 11612 30932 11664 30938
rect 11612 30874 11664 30880
rect 12440 30932 12492 30938
rect 12440 30874 12492 30880
rect 10876 30592 10928 30598
rect 10876 30534 10928 30540
rect 10600 30184 10652 30190
rect 10600 30126 10652 30132
rect 10612 29714 10640 30126
rect 10888 30054 10916 30534
rect 10968 30184 11020 30190
rect 10968 30126 11020 30132
rect 12440 30184 12492 30190
rect 12440 30126 12492 30132
rect 10876 30048 10928 30054
rect 10876 29990 10928 29996
rect 10600 29708 10652 29714
rect 10600 29650 10652 29656
rect 10692 29096 10744 29102
rect 10692 29038 10744 29044
rect 10704 28694 10732 29038
rect 10692 28688 10744 28694
rect 10692 28630 10744 28636
rect 10888 28626 10916 29990
rect 10980 29850 11008 30126
rect 11612 30116 11664 30122
rect 11612 30058 11664 30064
rect 10968 29844 11020 29850
rect 10968 29786 11020 29792
rect 11428 29776 11480 29782
rect 11428 29718 11480 29724
rect 10968 28960 11020 28966
rect 10968 28902 11020 28908
rect 10876 28620 10928 28626
rect 10876 28562 10928 28568
rect 10980 28014 11008 28902
rect 11060 28620 11112 28626
rect 11060 28562 11112 28568
rect 11072 28218 11100 28562
rect 11060 28212 11112 28218
rect 11060 28154 11112 28160
rect 10968 28008 11020 28014
rect 10968 27950 11020 27956
rect 11440 27606 11468 29718
rect 11624 29646 11652 30058
rect 12026 29948 12322 29968
rect 12082 29946 12106 29948
rect 12162 29946 12186 29948
rect 12242 29946 12266 29948
rect 12104 29894 12106 29946
rect 12168 29894 12180 29946
rect 12242 29894 12244 29946
rect 12082 29892 12106 29894
rect 12162 29892 12186 29894
rect 12242 29892 12266 29894
rect 12026 29872 12322 29892
rect 11612 29640 11664 29646
rect 11612 29582 11664 29588
rect 10416 27600 10468 27606
rect 10416 27542 10468 27548
rect 11428 27600 11480 27606
rect 11428 27542 11480 27548
rect 11244 27532 11296 27538
rect 11244 27474 11296 27480
rect 11520 27532 11572 27538
rect 11520 27474 11572 27480
rect 11060 27464 11112 27470
rect 11060 27406 11112 27412
rect 10600 26920 10652 26926
rect 10600 26862 10652 26868
rect 10324 26852 10376 26858
rect 10324 26794 10376 26800
rect 10232 26580 10284 26586
rect 10232 26522 10284 26528
rect 10140 26512 10192 26518
rect 10140 26454 10192 26460
rect 10612 26450 10640 26862
rect 10416 26444 10468 26450
rect 10416 26386 10468 26392
rect 10600 26444 10652 26450
rect 10600 26386 10652 26392
rect 10876 26444 10928 26450
rect 10876 26386 10928 26392
rect 9036 26240 9088 26246
rect 9036 26182 9088 26188
rect 9048 25906 9076 26182
rect 10428 26042 10456 26386
rect 10416 26036 10468 26042
rect 10416 25978 10468 25984
rect 9772 25968 9824 25974
rect 9772 25910 9824 25916
rect 9036 25900 9088 25906
rect 9036 25842 9088 25848
rect 9036 25696 9088 25702
rect 9036 25638 9088 25644
rect 9496 25696 9548 25702
rect 9496 25638 9548 25644
rect 9048 24410 9076 25638
rect 9508 25430 9536 25638
rect 9496 25424 9548 25430
rect 9416 25384 9496 25412
rect 9416 24682 9444 25384
rect 9496 25366 9548 25372
rect 9496 25152 9548 25158
rect 9496 25094 9548 25100
rect 9508 24750 9536 25094
rect 9784 24954 9812 25910
rect 10324 25832 10376 25838
rect 10324 25774 10376 25780
rect 9864 25356 9916 25362
rect 9864 25298 9916 25304
rect 9772 24948 9824 24954
rect 9772 24890 9824 24896
rect 9588 24880 9640 24886
rect 9588 24822 9640 24828
rect 9496 24744 9548 24750
rect 9496 24686 9548 24692
rect 9404 24676 9456 24682
rect 9404 24618 9456 24624
rect 9036 24404 9088 24410
rect 9036 24346 9088 24352
rect 9600 23866 9628 24822
rect 9876 24614 9904 25298
rect 10048 25220 10100 25226
rect 10048 25162 10100 25168
rect 9956 24676 10008 24682
rect 9956 24618 10008 24624
rect 9864 24608 9916 24614
rect 9864 24550 9916 24556
rect 9588 23860 9640 23866
rect 9588 23802 9640 23808
rect 9128 23724 9180 23730
rect 9128 23666 9180 23672
rect 9140 23322 9168 23666
rect 9220 23656 9272 23662
rect 9272 23604 9352 23610
rect 9220 23598 9352 23604
rect 9232 23582 9352 23598
rect 9128 23316 9180 23322
rect 9128 23258 9180 23264
rect 9324 23118 9352 23582
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 9324 22438 9352 23054
rect 9312 22432 9364 22438
rect 9312 22374 9364 22380
rect 9324 22166 9352 22374
rect 9312 22160 9364 22166
rect 9312 22102 9364 22108
rect 9324 21078 9352 22102
rect 9404 21480 9456 21486
rect 9404 21422 9456 21428
rect 9312 21072 9364 21078
rect 9312 21014 9364 21020
rect 8944 20324 8996 20330
rect 8944 20266 8996 20272
rect 8956 19310 8984 20266
rect 9324 19310 9352 21014
rect 9416 20466 9444 21422
rect 9600 21078 9628 23802
rect 9772 23656 9824 23662
rect 9772 23598 9824 23604
rect 9784 23254 9812 23598
rect 9772 23248 9824 23254
rect 9772 23190 9824 23196
rect 9680 21412 9732 21418
rect 9680 21354 9732 21360
rect 9588 21072 9640 21078
rect 9588 21014 9640 21020
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 9404 20460 9456 20466
rect 9404 20402 9456 20408
rect 9600 19310 9628 20878
rect 9692 20602 9720 21354
rect 9876 21350 9904 24550
rect 9968 24138 9996 24618
rect 9956 24132 10008 24138
rect 9956 24074 10008 24080
rect 9968 23662 9996 24074
rect 9956 23656 10008 23662
rect 9956 23598 10008 23604
rect 9956 23316 10008 23322
rect 9956 23258 10008 23264
rect 9864 21344 9916 21350
rect 9864 21286 9916 21292
rect 9876 21078 9904 21286
rect 9864 21072 9916 21078
rect 9864 21014 9916 21020
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9680 19984 9732 19990
rect 9680 19926 9732 19932
rect 8944 19304 8996 19310
rect 8944 19246 8996 19252
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9588 19304 9640 19310
rect 9588 19246 9640 19252
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 8404 17882 8432 19110
rect 8496 18834 8524 19110
rect 9692 18834 9720 19926
rect 9784 19922 9812 20878
rect 9968 20398 9996 23258
rect 10060 23186 10088 25162
rect 10232 24948 10284 24954
rect 10232 24890 10284 24896
rect 10244 24750 10272 24890
rect 10232 24744 10284 24750
rect 10232 24686 10284 24692
rect 10336 23730 10364 25774
rect 10784 25764 10836 25770
rect 10784 25706 10836 25712
rect 10796 24818 10824 25706
rect 10888 25362 10916 26386
rect 10876 25356 10928 25362
rect 10876 25298 10928 25304
rect 10784 24812 10836 24818
rect 10784 24754 10836 24760
rect 10600 24404 10652 24410
rect 10600 24346 10652 24352
rect 10612 23866 10640 24346
rect 10784 24336 10836 24342
rect 10784 24278 10836 24284
rect 10600 23860 10652 23866
rect 10600 23802 10652 23808
rect 10232 23724 10284 23730
rect 10232 23666 10284 23672
rect 10324 23724 10376 23730
rect 10324 23666 10376 23672
rect 10048 23180 10100 23186
rect 10048 23122 10100 23128
rect 10060 22094 10088 23122
rect 10244 22778 10272 23666
rect 10232 22772 10284 22778
rect 10232 22714 10284 22720
rect 10336 22234 10364 23666
rect 10324 22228 10376 22234
rect 10324 22170 10376 22176
rect 10796 22098 10824 24278
rect 10888 23050 10916 25298
rect 11072 23322 11100 27406
rect 11256 27062 11284 27474
rect 11532 27130 11560 27474
rect 11624 27470 11652 29582
rect 12452 29578 12480 30126
rect 12440 29572 12492 29578
rect 12440 29514 12492 29520
rect 12452 29306 12480 29514
rect 12440 29300 12492 29306
rect 12440 29242 12492 29248
rect 12544 29238 12572 31282
rect 12636 30802 12664 35226
rect 13372 35222 13400 36853
rect 15844 35488 15896 35494
rect 15844 35430 15896 35436
rect 13360 35216 13412 35222
rect 13360 35158 13412 35164
rect 13452 35216 13504 35222
rect 13452 35158 13504 35164
rect 12992 34536 13044 34542
rect 12992 34478 13044 34484
rect 12808 33992 12860 33998
rect 12808 33934 12860 33940
rect 12820 31754 12848 33934
rect 13004 32910 13032 34478
rect 13464 34202 13492 35158
rect 14464 35148 14516 35154
rect 14464 35090 14516 35096
rect 14280 35080 14332 35086
rect 14280 35022 14332 35028
rect 13820 34536 13872 34542
rect 13820 34478 13872 34484
rect 13452 34196 13504 34202
rect 13452 34138 13504 34144
rect 13832 34066 13860 34478
rect 13452 34060 13504 34066
rect 13452 34002 13504 34008
rect 13820 34060 13872 34066
rect 13820 34002 13872 34008
rect 13464 33454 13492 34002
rect 13544 33856 13596 33862
rect 13544 33798 13596 33804
rect 13556 33522 13584 33798
rect 13832 33522 13860 34002
rect 13544 33516 13596 33522
rect 13544 33458 13596 33464
rect 13820 33516 13872 33522
rect 13820 33458 13872 33464
rect 13268 33448 13320 33454
rect 13268 33390 13320 33396
rect 13452 33448 13504 33454
rect 13452 33390 13504 33396
rect 12900 32904 12952 32910
rect 12900 32846 12952 32852
rect 12992 32904 13044 32910
rect 12992 32846 13044 32852
rect 12912 32570 12940 32846
rect 12900 32564 12952 32570
rect 12900 32506 12952 32512
rect 13004 32314 13032 32846
rect 12912 32286 13032 32314
rect 13280 32298 13308 33390
rect 13544 32972 13596 32978
rect 13544 32914 13596 32920
rect 13556 32570 13584 32914
rect 14188 32768 14240 32774
rect 14188 32710 14240 32716
rect 13544 32564 13596 32570
rect 13544 32506 13596 32512
rect 13268 32292 13320 32298
rect 12808 31748 12860 31754
rect 12808 31690 12860 31696
rect 12624 30796 12676 30802
rect 12624 30738 12676 30744
rect 12808 30048 12860 30054
rect 12808 29990 12860 29996
rect 12716 29776 12768 29782
rect 12716 29718 12768 29724
rect 12728 29306 12756 29718
rect 12716 29300 12768 29306
rect 12716 29242 12768 29248
rect 11888 29232 11940 29238
rect 11888 29174 11940 29180
rect 12532 29232 12584 29238
rect 12532 29174 12584 29180
rect 11704 27532 11756 27538
rect 11704 27474 11756 27480
rect 11612 27464 11664 27470
rect 11612 27406 11664 27412
rect 11520 27124 11572 27130
rect 11520 27066 11572 27072
rect 11244 27056 11296 27062
rect 11244 26998 11296 27004
rect 11152 26920 11204 26926
rect 11152 26862 11204 26868
rect 11164 25974 11192 26862
rect 11256 26382 11284 26998
rect 11244 26376 11296 26382
rect 11244 26318 11296 26324
rect 11428 26376 11480 26382
rect 11428 26318 11480 26324
rect 11440 25974 11468 26318
rect 11152 25968 11204 25974
rect 11152 25910 11204 25916
rect 11428 25968 11480 25974
rect 11428 25910 11480 25916
rect 11164 25401 11192 25910
rect 11150 25392 11206 25401
rect 11440 25362 11468 25910
rect 11716 25838 11744 27474
rect 11900 26246 11928 29174
rect 12716 29028 12768 29034
rect 12716 28970 12768 28976
rect 12026 28860 12322 28880
rect 12082 28858 12106 28860
rect 12162 28858 12186 28860
rect 12242 28858 12266 28860
rect 12104 28806 12106 28858
rect 12168 28806 12180 28858
rect 12242 28806 12244 28858
rect 12082 28804 12106 28806
rect 12162 28804 12186 28806
rect 12242 28804 12266 28806
rect 12026 28784 12322 28804
rect 12624 28416 12676 28422
rect 12624 28358 12676 28364
rect 12636 28014 12664 28358
rect 12624 28008 12676 28014
rect 12624 27950 12676 27956
rect 12348 27940 12400 27946
rect 12348 27882 12400 27888
rect 12026 27772 12322 27792
rect 12082 27770 12106 27772
rect 12162 27770 12186 27772
rect 12242 27770 12266 27772
rect 12104 27718 12106 27770
rect 12168 27718 12180 27770
rect 12242 27718 12244 27770
rect 12082 27716 12106 27718
rect 12162 27716 12186 27718
rect 12242 27716 12266 27718
rect 12026 27696 12322 27716
rect 12360 27334 12388 27882
rect 12440 27532 12492 27538
rect 12440 27474 12492 27480
rect 12072 27328 12124 27334
rect 12072 27270 12124 27276
rect 12348 27328 12400 27334
rect 12348 27270 12400 27276
rect 12084 26858 12112 27270
rect 12348 27124 12400 27130
rect 12348 27066 12400 27072
rect 12072 26852 12124 26858
rect 12072 26794 12124 26800
rect 12026 26684 12322 26704
rect 12082 26682 12106 26684
rect 12162 26682 12186 26684
rect 12242 26682 12266 26684
rect 12104 26630 12106 26682
rect 12168 26630 12180 26682
rect 12242 26630 12244 26682
rect 12082 26628 12106 26630
rect 12162 26628 12186 26630
rect 12242 26628 12266 26630
rect 12026 26608 12322 26628
rect 12164 26512 12216 26518
rect 12084 26460 12164 26466
rect 12084 26454 12216 26460
rect 11980 26444 12032 26450
rect 12084 26438 12204 26454
rect 12084 26432 12112 26438
rect 12032 26404 12112 26432
rect 11980 26386 12032 26392
rect 11888 26240 11940 26246
rect 11888 26182 11940 26188
rect 11704 25832 11756 25838
rect 11704 25774 11756 25780
rect 11150 25327 11152 25336
rect 11204 25327 11206 25336
rect 11428 25356 11480 25362
rect 11152 25298 11204 25304
rect 11428 25298 11480 25304
rect 11716 24970 11744 25774
rect 11796 25764 11848 25770
rect 11796 25706 11848 25712
rect 11624 24942 11744 24970
rect 11244 24608 11296 24614
rect 11244 24550 11296 24556
rect 11256 24342 11284 24550
rect 11624 24410 11652 24942
rect 11612 24404 11664 24410
rect 11612 24346 11664 24352
rect 11244 24336 11296 24342
rect 11244 24278 11296 24284
rect 11244 24200 11296 24206
rect 11244 24142 11296 24148
rect 11520 24200 11572 24206
rect 11520 24142 11572 24148
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 11256 23186 11284 24142
rect 11532 23798 11560 24142
rect 11624 24070 11652 24346
rect 11808 24274 11836 25706
rect 11900 25702 11928 26182
rect 12360 25838 12388 27066
rect 12452 26926 12480 27474
rect 12440 26920 12492 26926
rect 12440 26862 12492 26868
rect 12440 26512 12492 26518
rect 12440 26454 12492 26460
rect 12452 25974 12480 26454
rect 12624 26240 12676 26246
rect 12624 26182 12676 26188
rect 12440 25968 12492 25974
rect 12440 25910 12492 25916
rect 12348 25832 12400 25838
rect 12636 25786 12664 26182
rect 12348 25774 12400 25780
rect 12544 25758 12664 25786
rect 11888 25696 11940 25702
rect 11888 25638 11940 25644
rect 12026 25596 12322 25616
rect 12082 25594 12106 25596
rect 12162 25594 12186 25596
rect 12242 25594 12266 25596
rect 12104 25542 12106 25594
rect 12168 25542 12180 25594
rect 12242 25542 12244 25594
rect 12082 25540 12106 25542
rect 12162 25540 12186 25542
rect 12242 25540 12266 25542
rect 12026 25520 12322 25540
rect 12544 25362 12572 25758
rect 12624 25492 12676 25498
rect 12624 25434 12676 25440
rect 12440 25356 12492 25362
rect 12440 25298 12492 25304
rect 12532 25356 12584 25362
rect 12532 25298 12584 25304
rect 12164 25220 12216 25226
rect 12164 25162 12216 25168
rect 12176 24886 12204 25162
rect 12164 24880 12216 24886
rect 12164 24822 12216 24828
rect 11888 24812 11940 24818
rect 11888 24754 11940 24760
rect 11796 24268 11848 24274
rect 11796 24210 11848 24216
rect 11704 24132 11756 24138
rect 11704 24074 11756 24080
rect 11612 24064 11664 24070
rect 11612 24006 11664 24012
rect 11716 23866 11744 24074
rect 11704 23860 11756 23866
rect 11704 23802 11756 23808
rect 11520 23792 11572 23798
rect 11520 23734 11572 23740
rect 11428 23656 11480 23662
rect 11428 23598 11480 23604
rect 11440 23254 11468 23598
rect 11900 23322 11928 24754
rect 12256 24744 12308 24750
rect 12308 24692 12388 24698
rect 12256 24686 12388 24692
rect 12268 24670 12388 24686
rect 12026 24508 12322 24528
rect 12082 24506 12106 24508
rect 12162 24506 12186 24508
rect 12242 24506 12266 24508
rect 12104 24454 12106 24506
rect 12168 24454 12180 24506
rect 12242 24454 12244 24506
rect 12082 24452 12106 24454
rect 12162 24452 12186 24454
rect 12242 24452 12266 24454
rect 12026 24432 12322 24452
rect 12360 24290 12388 24670
rect 12268 24262 12388 24290
rect 12268 24070 12296 24262
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12256 24064 12308 24070
rect 12256 24006 12308 24012
rect 12268 23610 12296 24006
rect 12360 23866 12388 24142
rect 12348 23860 12400 23866
rect 12452 23848 12480 25298
rect 12452 23820 12572 23848
rect 12348 23802 12400 23808
rect 12440 23724 12492 23730
rect 12440 23666 12492 23672
rect 12268 23582 12388 23610
rect 12026 23420 12322 23440
rect 12082 23418 12106 23420
rect 12162 23418 12186 23420
rect 12242 23418 12266 23420
rect 12104 23366 12106 23418
rect 12168 23366 12180 23418
rect 12242 23366 12244 23418
rect 12082 23364 12106 23366
rect 12162 23364 12186 23366
rect 12242 23364 12266 23366
rect 12026 23344 12322 23364
rect 11888 23316 11940 23322
rect 11888 23258 11940 23264
rect 11428 23248 11480 23254
rect 11428 23190 11480 23196
rect 11244 23180 11296 23186
rect 11244 23122 11296 23128
rect 10876 23044 10928 23050
rect 10876 22986 10928 22992
rect 10968 22772 11020 22778
rect 10968 22714 11020 22720
rect 10980 22506 11008 22714
rect 11152 22568 11204 22574
rect 11152 22510 11204 22516
rect 10968 22500 11020 22506
rect 10968 22442 11020 22448
rect 10876 22228 10928 22234
rect 10876 22170 10928 22176
rect 10060 22066 10272 22094
rect 10140 21548 10192 21554
rect 10140 21490 10192 21496
rect 9956 20392 10008 20398
rect 9956 20334 10008 20340
rect 10152 19922 10180 21490
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 10140 19916 10192 19922
rect 10140 19858 10192 19864
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 9864 19236 9916 19242
rect 9864 19178 9916 19184
rect 9876 18970 9904 19178
rect 10060 18970 10088 19246
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 8484 18828 8536 18834
rect 8484 18770 8536 18776
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9600 18222 9628 18362
rect 9876 18290 9904 18906
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 5908 17740 5960 17746
rect 5908 17682 5960 17688
rect 6184 17740 6236 17746
rect 6184 17682 6236 17688
rect 6368 17740 6420 17746
rect 6368 17682 6420 17688
rect 7472 17740 7524 17746
rect 7472 17682 7524 17688
rect 5920 17338 5948 17682
rect 7196 17604 7248 17610
rect 7196 17546 7248 17552
rect 6491 17436 6787 17456
rect 6547 17434 6571 17436
rect 6627 17434 6651 17436
rect 6707 17434 6731 17436
rect 6569 17382 6571 17434
rect 6633 17382 6645 17434
rect 6707 17382 6709 17434
rect 6547 17380 6571 17382
rect 6627 17380 6651 17382
rect 6707 17380 6731 17382
rect 6491 17360 6787 17380
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 7208 17134 7236 17546
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7392 17202 7420 17478
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 5644 16658 5672 17070
rect 6368 17060 6420 17066
rect 6368 17002 6420 17008
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 6380 16590 6408 17002
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 6840 16726 6868 16934
rect 7300 16794 7328 16934
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 6828 16720 6880 16726
rect 6828 16662 6880 16668
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6380 16046 6408 16526
rect 6491 16348 6787 16368
rect 6547 16346 6571 16348
rect 6627 16346 6651 16348
rect 6707 16346 6731 16348
rect 6569 16294 6571 16346
rect 6633 16294 6645 16346
rect 6707 16294 6709 16346
rect 6547 16292 6571 16294
rect 6627 16292 6651 16294
rect 6707 16292 6731 16294
rect 6491 16272 6787 16292
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 6368 16040 6420 16046
rect 6368 15982 6420 15988
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 5184 15366 5212 15982
rect 6656 15502 6684 15982
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 6368 15496 6420 15502
rect 6368 15438 6420 15444
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 5080 15020 5132 15026
rect 5080 14962 5132 14968
rect 5092 14482 5120 14962
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 5184 14618 5212 14894
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 5460 14550 5488 14758
rect 5448 14544 5500 14550
rect 5448 14486 5500 14492
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 6012 13870 6040 15302
rect 6380 14346 6408 15438
rect 6491 15260 6787 15280
rect 6547 15258 6571 15260
rect 6627 15258 6651 15260
rect 6707 15258 6731 15260
rect 6569 15206 6571 15258
rect 6633 15206 6645 15258
rect 6707 15206 6709 15258
rect 6547 15204 6571 15206
rect 6627 15204 6651 15206
rect 6707 15204 6731 15206
rect 6491 15184 6787 15204
rect 6368 14340 6420 14346
rect 6368 14282 6420 14288
rect 6491 14172 6787 14192
rect 6547 14170 6571 14172
rect 6627 14170 6651 14172
rect 6707 14170 6731 14172
rect 6569 14118 6571 14170
rect 6633 14118 6645 14170
rect 6707 14118 6709 14170
rect 6547 14116 6571 14118
rect 6627 14116 6651 14118
rect 6707 14116 6731 14118
rect 6491 14096 6787 14116
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4988 13728 5040 13734
rect 4988 13670 5040 13676
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 4080 12782 4108 13670
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4724 12850 4752 13262
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 3884 12368 3936 12374
rect 3884 12310 3936 12316
rect 4080 12306 4108 12718
rect 5368 12714 5396 13670
rect 5460 12986 5488 13806
rect 6012 13326 6040 13806
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6932 13326 6960 13670
rect 7024 13462 7052 15642
rect 7484 15638 7512 17682
rect 8404 17066 8432 17818
rect 8496 17202 8524 18022
rect 9600 17542 9628 18158
rect 10048 18148 10100 18154
rect 10048 18090 10100 18096
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8392 17060 8444 17066
rect 8392 17002 8444 17008
rect 7564 15972 7616 15978
rect 7564 15914 7616 15920
rect 8024 15972 8076 15978
rect 8024 15914 8076 15920
rect 8852 15972 8904 15978
rect 8852 15914 8904 15920
rect 7288 15632 7340 15638
rect 7288 15574 7340 15580
rect 7472 15632 7524 15638
rect 7472 15574 7524 15580
rect 7300 14822 7328 15574
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7300 14618 7328 14758
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7484 14482 7512 15302
rect 7576 14618 7604 15914
rect 8036 15706 8064 15914
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 8220 15570 8248 15846
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7852 14958 7880 15438
rect 8220 14958 8248 15506
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7852 13870 7880 14894
rect 8312 14550 8340 15370
rect 8300 14544 8352 14550
rect 8300 14486 8352 14492
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 7852 13530 7880 13806
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 7024 13326 7052 13398
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 6012 12714 6040 13262
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 6491 13084 6787 13104
rect 6547 13082 6571 13084
rect 6627 13082 6651 13084
rect 6707 13082 6731 13084
rect 6569 13030 6571 13082
rect 6633 13030 6645 13082
rect 6707 13030 6709 13082
rect 6547 13028 6571 13030
rect 6627 13028 6651 13030
rect 6707 13028 6731 13030
rect 6491 13008 6787 13028
rect 7852 12782 7880 13126
rect 7944 12850 7972 13806
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 5368 12374 5396 12650
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 3988 10674 4016 12174
rect 5000 11898 5028 12174
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 5184 11150 5212 11630
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4908 10674 4936 10950
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 5276 9586 5304 11154
rect 5368 10538 5396 12310
rect 5460 12102 5488 12582
rect 6012 12238 6040 12650
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5460 11762 5488 12038
rect 6012 11762 6040 12174
rect 6491 11996 6787 12016
rect 6547 11994 6571 11996
rect 6627 11994 6651 11996
rect 6707 11994 6731 11996
rect 6569 11942 6571 11994
rect 6633 11942 6645 11994
rect 6707 11942 6709 11994
rect 6547 11940 6571 11942
rect 6627 11940 6651 11942
rect 6707 11940 6731 11942
rect 6491 11920 6787 11940
rect 7116 11762 7144 12582
rect 7944 12442 7972 12786
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 5540 11620 5592 11626
rect 5540 11562 5592 11568
rect 5552 11218 5580 11562
rect 8036 11558 8064 13262
rect 8680 12986 8708 13330
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8772 12782 8800 13670
rect 8864 13258 8892 15914
rect 9692 15638 9720 17818
rect 9968 17338 9996 18022
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 10060 16726 10088 18090
rect 10048 16720 10100 16726
rect 10048 16662 10100 16668
rect 10152 16114 10180 19858
rect 10244 18766 10272 22066
rect 10784 22092 10836 22098
rect 10784 22034 10836 22040
rect 10796 21486 10824 22034
rect 10784 21480 10836 21486
rect 10784 21422 10836 21428
rect 10508 20800 10560 20806
rect 10508 20742 10560 20748
rect 10520 20398 10548 20742
rect 10508 20392 10560 20398
rect 10508 20334 10560 20340
rect 10520 19514 10548 20334
rect 10692 19916 10744 19922
rect 10692 19858 10744 19864
rect 10508 19508 10560 19514
rect 10508 19450 10560 19456
rect 10704 19446 10732 19858
rect 10692 19440 10744 19446
rect 10692 19382 10744 19388
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10336 18822 10640 18850
rect 10704 18834 10732 19110
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10336 18698 10364 18822
rect 10612 18766 10640 18822
rect 10692 18828 10744 18834
rect 10692 18770 10744 18776
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10324 18692 10376 18698
rect 10324 18634 10376 18640
rect 10416 18692 10468 18698
rect 10416 18634 10468 18640
rect 10428 17746 10456 18634
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10704 18426 10732 18566
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 10416 17740 10468 17746
rect 10416 17682 10468 17688
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9680 15632 9732 15638
rect 9680 15574 9732 15580
rect 9784 14890 9812 15642
rect 10508 15360 10560 15366
rect 10508 15302 10560 15308
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 9772 14884 9824 14890
rect 9772 14826 9824 14832
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 8852 13252 8904 13258
rect 8852 13194 8904 13200
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8864 12434 8892 13194
rect 9140 12850 9168 13670
rect 9600 12918 9628 13670
rect 9956 13320 10008 13326
rect 10060 13274 10088 15098
rect 10520 15026 10548 15302
rect 10796 15026 10824 17614
rect 10888 16046 10916 22170
rect 10980 21010 11008 22442
rect 11060 22160 11112 22166
rect 11060 22102 11112 22108
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 11072 20398 11100 22102
rect 11164 22098 11192 22510
rect 11152 22092 11204 22098
rect 11152 22034 11204 22040
rect 11164 21690 11192 22034
rect 11244 21888 11296 21894
rect 11244 21830 11296 21836
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 11256 21554 11284 21830
rect 11244 21548 11296 21554
rect 11244 21490 11296 21496
rect 11440 21146 11468 23190
rect 11796 22432 11848 22438
rect 11796 22374 11848 22380
rect 11704 22228 11756 22234
rect 11704 22170 11756 22176
rect 11716 21622 11744 22170
rect 11704 21616 11756 21622
rect 11704 21558 11756 21564
rect 11808 21486 11836 22374
rect 12026 22332 12322 22352
rect 12082 22330 12106 22332
rect 12162 22330 12186 22332
rect 12242 22330 12266 22332
rect 12104 22278 12106 22330
rect 12168 22278 12180 22330
rect 12242 22278 12244 22330
rect 12082 22276 12106 22278
rect 12162 22276 12186 22278
rect 12242 22276 12266 22278
rect 12026 22256 12322 22276
rect 12360 22234 12388 23582
rect 12452 23254 12480 23666
rect 12440 23248 12492 23254
rect 12440 23190 12492 23196
rect 12348 22228 12400 22234
rect 12348 22170 12400 22176
rect 12348 22092 12400 22098
rect 12348 22034 12400 22040
rect 11888 22024 11940 22030
rect 11888 21966 11940 21972
rect 12162 21992 12218 22001
rect 11796 21480 11848 21486
rect 11796 21422 11848 21428
rect 11428 21140 11480 21146
rect 11428 21082 11480 21088
rect 11808 20992 11836 21422
rect 11900 21146 11928 21966
rect 12162 21927 12164 21936
rect 12216 21927 12218 21936
rect 12164 21898 12216 21904
rect 12026 21244 12322 21264
rect 12082 21242 12106 21244
rect 12162 21242 12186 21244
rect 12242 21242 12266 21244
rect 12104 21190 12106 21242
rect 12168 21190 12180 21242
rect 12242 21190 12244 21242
rect 12082 21188 12106 21190
rect 12162 21188 12186 21190
rect 12242 21188 12266 21190
rect 12026 21168 12322 21188
rect 11888 21140 11940 21146
rect 11888 21082 11940 21088
rect 11888 21004 11940 21010
rect 11808 20964 11888 20992
rect 11888 20946 11940 20952
rect 11900 20602 11928 20946
rect 12256 20936 12308 20942
rect 12360 20924 12388 22034
rect 12452 21690 12480 23190
rect 12544 22710 12572 23820
rect 12636 23594 12664 25434
rect 12624 23588 12676 23594
rect 12624 23530 12676 23536
rect 12636 23168 12664 23530
rect 12728 23338 12756 28970
rect 12820 28626 12848 29990
rect 12912 29646 12940 32286
rect 13268 32234 13320 32240
rect 12992 32224 13044 32230
rect 12992 32166 13044 32172
rect 13176 32224 13228 32230
rect 13176 32166 13228 32172
rect 13004 32026 13032 32166
rect 12992 32020 13044 32026
rect 12992 31962 13044 31968
rect 13188 31754 13216 32166
rect 13280 31754 13308 32234
rect 13176 31748 13228 31754
rect 13280 31726 13400 31754
rect 13176 31690 13228 31696
rect 13084 31136 13136 31142
rect 13084 31078 13136 31084
rect 12992 30184 13044 30190
rect 12992 30126 13044 30132
rect 13004 30054 13032 30126
rect 12992 30048 13044 30054
rect 12992 29990 13044 29996
rect 13096 29850 13124 31078
rect 13084 29844 13136 29850
rect 13084 29786 13136 29792
rect 12900 29640 12952 29646
rect 12900 29582 12952 29588
rect 12912 29510 12940 29582
rect 12900 29504 12952 29510
rect 12900 29446 12952 29452
rect 13096 29102 13124 29786
rect 13188 29170 13216 31690
rect 13372 31278 13400 31726
rect 13360 31272 13412 31278
rect 13360 31214 13412 31220
rect 13912 31272 13964 31278
rect 13912 31214 13964 31220
rect 13372 30734 13400 31214
rect 13924 30938 13952 31214
rect 13912 30932 13964 30938
rect 13912 30874 13964 30880
rect 13636 30796 13688 30802
rect 13636 30738 13688 30744
rect 13360 30728 13412 30734
rect 13360 30670 13412 30676
rect 13176 29164 13228 29170
rect 13176 29106 13228 29112
rect 12900 29096 12952 29102
rect 12900 29038 12952 29044
rect 13084 29096 13136 29102
rect 13084 29038 13136 29044
rect 12808 28620 12860 28626
rect 12808 28562 12860 28568
rect 12912 26926 12940 29038
rect 12992 28620 13044 28626
rect 12992 28562 13044 28568
rect 13004 27674 13032 28562
rect 13372 28490 13400 30670
rect 13648 28626 13676 30738
rect 14200 30190 14228 32710
rect 14188 30184 14240 30190
rect 14188 30126 14240 30132
rect 13912 30116 13964 30122
rect 13912 30058 13964 30064
rect 13728 29504 13780 29510
rect 13728 29446 13780 29452
rect 13636 28620 13688 28626
rect 13636 28562 13688 28568
rect 13360 28484 13412 28490
rect 13360 28426 13412 28432
rect 13084 28008 13136 28014
rect 13084 27950 13136 27956
rect 12992 27668 13044 27674
rect 12992 27610 13044 27616
rect 13096 27062 13124 27950
rect 13084 27056 13136 27062
rect 13084 26998 13136 27004
rect 12900 26920 12952 26926
rect 12900 26862 12952 26868
rect 13268 26920 13320 26926
rect 13268 26862 13320 26868
rect 12808 26308 12860 26314
rect 12808 26250 12860 26256
rect 12820 25430 12848 26250
rect 13176 25764 13228 25770
rect 13176 25706 13228 25712
rect 12900 25696 12952 25702
rect 12900 25638 12952 25644
rect 12808 25424 12860 25430
rect 12806 25392 12808 25401
rect 12860 25392 12862 25401
rect 12912 25362 12940 25638
rect 13188 25498 13216 25706
rect 13176 25492 13228 25498
rect 13176 25434 13228 25440
rect 12806 25327 12862 25336
rect 12900 25356 12952 25362
rect 12900 25298 12952 25304
rect 12992 24744 13044 24750
rect 12992 24686 13044 24692
rect 13004 24410 13032 24686
rect 12992 24404 13044 24410
rect 12992 24346 13044 24352
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 12912 23730 12940 24006
rect 12900 23724 12952 23730
rect 12900 23666 12952 23672
rect 13280 23526 13308 26862
rect 13372 24682 13400 28426
rect 13740 28082 13768 29446
rect 13924 28218 13952 30058
rect 14004 28620 14056 28626
rect 14004 28562 14056 28568
rect 13912 28212 13964 28218
rect 13912 28154 13964 28160
rect 13728 28076 13780 28082
rect 13728 28018 13780 28024
rect 13452 27532 13504 27538
rect 13452 27474 13504 27480
rect 13464 27130 13492 27474
rect 13452 27124 13504 27130
rect 13452 27066 13504 27072
rect 13544 27124 13596 27130
rect 13544 27066 13596 27072
rect 13556 27010 13584 27066
rect 13464 26994 13584 27010
rect 13452 26988 13584 26994
rect 13504 26982 13584 26988
rect 13452 26930 13504 26936
rect 13636 26784 13688 26790
rect 13636 26726 13688 26732
rect 13648 25906 13676 26726
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 13648 24750 13676 25842
rect 13740 25226 13768 28018
rect 13820 26920 13872 26926
rect 13820 26862 13872 26868
rect 13832 26518 13860 26862
rect 13820 26512 13872 26518
rect 13820 26454 13872 26460
rect 13820 26036 13872 26042
rect 13820 25978 13872 25984
rect 13832 25294 13860 25978
rect 13820 25288 13872 25294
rect 13820 25230 13872 25236
rect 13728 25220 13780 25226
rect 13728 25162 13780 25168
rect 13636 24744 13688 24750
rect 13636 24686 13688 24692
rect 13360 24676 13412 24682
rect 13360 24618 13412 24624
rect 13832 24614 13860 25230
rect 14016 24886 14044 28562
rect 14188 27872 14240 27878
rect 14188 27814 14240 27820
rect 14200 27606 14228 27814
rect 14188 27600 14240 27606
rect 14188 27542 14240 27548
rect 14188 26988 14240 26994
rect 14188 26930 14240 26936
rect 14004 24880 14056 24886
rect 14004 24822 14056 24828
rect 13820 24608 13872 24614
rect 13820 24550 13872 24556
rect 13832 23610 13860 24550
rect 13740 23594 13860 23610
rect 13728 23588 13860 23594
rect 13780 23582 13860 23588
rect 13728 23530 13780 23536
rect 13268 23520 13320 23526
rect 13268 23462 13320 23468
rect 13636 23520 13688 23526
rect 13636 23462 13688 23468
rect 12728 23310 12848 23338
rect 12716 23180 12768 23186
rect 12636 23140 12716 23168
rect 12716 23122 12768 23128
rect 12532 22704 12584 22710
rect 12532 22646 12584 22652
rect 12820 22094 12848 23310
rect 12992 22976 13044 22982
rect 12992 22918 13044 22924
rect 13004 22778 13032 22918
rect 12992 22772 13044 22778
rect 12992 22714 13044 22720
rect 13176 22636 13228 22642
rect 13176 22578 13228 22584
rect 12636 22066 12848 22094
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 12544 21622 12572 21966
rect 12532 21616 12584 21622
rect 12532 21558 12584 21564
rect 12532 21480 12584 21486
rect 12532 21422 12584 21428
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12452 20942 12480 21286
rect 12544 21010 12572 21422
rect 12532 21004 12584 21010
rect 12532 20946 12584 20952
rect 12308 20896 12388 20924
rect 12256 20878 12308 20884
rect 12360 20602 12388 20896
rect 12440 20936 12492 20942
rect 12440 20878 12492 20884
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 11060 20392 11112 20398
rect 11060 20334 11112 20340
rect 11336 20392 11388 20398
rect 11336 20334 11388 20340
rect 10968 20324 11020 20330
rect 10968 20266 11020 20272
rect 10980 20210 11008 20266
rect 10980 20182 11100 20210
rect 10968 18896 11020 18902
rect 10968 18838 11020 18844
rect 10980 18426 11008 18838
rect 10968 18420 11020 18426
rect 10968 18362 11020 18368
rect 11072 18086 11100 20182
rect 11348 18834 11376 20334
rect 12452 20330 12480 20878
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12440 20324 12492 20330
rect 12440 20266 12492 20272
rect 12026 20156 12322 20176
rect 12082 20154 12106 20156
rect 12162 20154 12186 20156
rect 12242 20154 12266 20156
rect 12104 20102 12106 20154
rect 12168 20102 12180 20154
rect 12242 20102 12244 20154
rect 12082 20100 12106 20102
rect 12162 20100 12186 20102
rect 12242 20100 12266 20102
rect 12026 20080 12322 20100
rect 12544 19990 12572 20334
rect 12532 19984 12584 19990
rect 12532 19926 12584 19932
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 11796 19848 11848 19854
rect 11796 19790 11848 19796
rect 11808 19310 11836 19790
rect 12268 19514 12296 19858
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 11796 19304 11848 19310
rect 11796 19246 11848 19252
rect 11520 19236 11572 19242
rect 11520 19178 11572 19184
rect 11532 18834 11560 19178
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 11152 18216 11204 18222
rect 11152 18158 11204 18164
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10888 15570 10916 15846
rect 10968 15632 11020 15638
rect 10968 15574 11020 15580
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10796 13326 10824 14962
rect 10980 13410 11008 15574
rect 11072 15094 11100 18022
rect 11164 17338 11192 18158
rect 11612 17604 11664 17610
rect 11612 17546 11664 17552
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11532 16658 11560 17478
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11336 16176 11388 16182
rect 11336 16118 11388 16124
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 11256 14822 11284 15506
rect 11348 15502 11376 16118
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 10980 13382 11192 13410
rect 10980 13326 11008 13382
rect 10008 13268 10088 13274
rect 9956 13262 10088 13268
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 9968 13246 10088 13262
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 8772 12406 8892 12434
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8496 11694 8524 12038
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5552 10810 5580 11154
rect 6491 10908 6787 10928
rect 6547 10906 6571 10908
rect 6627 10906 6651 10908
rect 6707 10906 6731 10908
rect 6569 10854 6571 10906
rect 6633 10854 6645 10906
rect 6707 10854 6709 10906
rect 6547 10852 6571 10854
rect 6627 10852 6651 10854
rect 6707 10852 6731 10854
rect 6491 10832 6787 10852
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 3332 9444 3384 9450
rect 3332 9386 3384 9392
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3160 8430 3188 8774
rect 3344 8498 3372 9386
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 2320 8016 2372 8022
rect 2320 7958 2372 7964
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 1504 6914 1532 7890
rect 1860 7200 1912 7206
rect 1860 7142 1912 7148
rect 1412 6886 1532 6914
rect 1412 6798 1440 6886
rect 1872 6866 1900 7142
rect 2332 7002 2360 7958
rect 2792 7886 2820 8230
rect 3252 8090 3280 8230
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 5234 1440 6734
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2608 5234 2636 5510
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 1412 4146 1440 5170
rect 2700 5166 2728 6938
rect 2976 6662 3004 7278
rect 3160 7018 3188 7346
rect 3252 7206 3280 8026
rect 3344 7410 3372 8434
rect 3804 8430 3832 9454
rect 4448 8634 4476 9454
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4632 9042 4660 9318
rect 5276 9178 5304 9522
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5368 9110 5396 10474
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 6491 9820 6787 9840
rect 6547 9818 6571 9820
rect 6627 9818 6651 9820
rect 6707 9818 6731 9820
rect 6569 9766 6571 9818
rect 6633 9766 6645 9818
rect 6707 9766 6709 9818
rect 6547 9764 6571 9766
rect 6627 9764 6651 9766
rect 6707 9764 6731 9766
rect 6491 9744 6787 9764
rect 7116 9586 7144 9862
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 4448 7478 4476 8570
rect 4540 8566 4568 8910
rect 4528 8560 4580 8566
rect 4528 8502 4580 8508
rect 4540 7954 4568 8502
rect 5368 8090 5396 9046
rect 5644 8090 5672 9386
rect 6491 8732 6787 8752
rect 6547 8730 6571 8732
rect 6627 8730 6651 8732
rect 6707 8730 6731 8732
rect 6569 8678 6571 8730
rect 6633 8678 6645 8730
rect 6707 8678 6709 8730
rect 6547 8676 6571 8678
rect 6627 8676 6651 8678
rect 6707 8676 6731 8678
rect 6491 8656 6787 8676
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4436 7472 4488 7478
rect 4436 7414 4488 7420
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3160 6990 3280 7018
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2976 5914 3004 6598
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 3252 5710 3280 6990
rect 4540 6730 4568 7890
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5184 7546 5212 7822
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5368 7256 5396 8026
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 5276 7228 5396 7256
rect 4528 6724 4580 6730
rect 4528 6666 4580 6672
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4264 6322 4292 6598
rect 4540 6322 4568 6666
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 3068 5370 3096 5646
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 3068 4758 3096 5306
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 3252 4622 3280 5646
rect 4540 4690 4568 6258
rect 5276 6186 5304 7228
rect 5460 6798 5488 7414
rect 5644 7410 5672 8026
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5552 6866 5580 7142
rect 5632 6928 5684 6934
rect 5632 6870 5684 6876
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5264 6180 5316 6186
rect 5264 6122 5316 6128
rect 5276 5846 5304 6122
rect 5264 5840 5316 5846
rect 5184 5788 5264 5794
rect 5184 5782 5316 5788
rect 5184 5766 5304 5782
rect 5184 5098 5212 5766
rect 5356 5228 5408 5234
rect 5460 5216 5488 6734
rect 5552 6458 5580 6802
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5644 5914 5672 6870
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5644 5234 5672 5850
rect 5408 5188 5488 5216
rect 5632 5228 5684 5234
rect 5356 5170 5408 5176
rect 5632 5170 5684 5176
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 5184 4758 5212 5034
rect 5172 4752 5224 4758
rect 5172 4694 5224 4700
rect 4528 4684 4580 4690
rect 4528 4626 4580 4632
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 1872 4185 1900 4422
rect 1858 4176 1914 4185
rect 1400 4140 1452 4146
rect 2608 4146 2636 4422
rect 3068 4282 3096 4558
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 1858 4111 1914 4120
rect 2596 4140 2648 4146
rect 1400 4082 1452 4088
rect 2596 4082 2648 4088
rect 4080 3602 4108 4218
rect 4632 3738 4660 4558
rect 5184 4010 5212 4694
rect 5368 4146 5396 5170
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5552 4146 5580 4966
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 5184 3670 5212 3946
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 5368 3534 5396 4082
rect 5552 3738 5580 4082
rect 5644 4010 5672 4422
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5644 3602 5672 3946
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5736 2650 5764 8570
rect 6840 8566 6868 9454
rect 8036 9432 8064 11494
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8220 10130 8248 10406
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8116 10056 8168 10062
rect 8312 10010 8340 10542
rect 8576 10532 8628 10538
rect 8576 10474 8628 10480
rect 8168 10004 8340 10010
rect 8116 9998 8340 10004
rect 8128 9982 8340 9998
rect 8116 9444 8168 9450
rect 8036 9404 8116 9432
rect 8116 9386 8168 9392
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6491 7644 6787 7664
rect 6547 7642 6571 7644
rect 6627 7642 6651 7644
rect 6707 7642 6731 7644
rect 6569 7590 6571 7642
rect 6633 7590 6645 7642
rect 6707 7590 6709 7642
rect 6547 7588 6571 7590
rect 6627 7588 6651 7590
rect 6707 7588 6731 7590
rect 6491 7568 6787 7588
rect 6840 6882 6868 8502
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7576 7342 7604 7686
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 6840 6854 6960 6882
rect 6491 6556 6787 6576
rect 6547 6554 6571 6556
rect 6627 6554 6651 6556
rect 6707 6554 6731 6556
rect 6569 6502 6571 6554
rect 6633 6502 6645 6554
rect 6707 6502 6709 6554
rect 6547 6500 6571 6502
rect 6627 6500 6651 6502
rect 6707 6500 6731 6502
rect 6491 6480 6787 6500
rect 6932 6322 6960 6854
rect 7208 6322 7236 7142
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 6491 5468 6787 5488
rect 6547 5466 6571 5468
rect 6627 5466 6651 5468
rect 6707 5466 6731 5468
rect 6569 5414 6571 5466
rect 6633 5414 6645 5466
rect 6707 5414 6709 5466
rect 6547 5412 6571 5414
rect 6627 5412 6651 5414
rect 6707 5412 6731 5414
rect 6491 5392 6787 5412
rect 6491 4380 6787 4400
rect 6547 4378 6571 4380
rect 6627 4378 6651 4380
rect 6707 4378 6731 4380
rect 6569 4326 6571 4378
rect 6633 4326 6645 4378
rect 6707 4326 6709 4378
rect 6547 4324 6571 4326
rect 6627 4324 6651 4326
rect 6707 4324 6731 4326
rect 6491 4304 6787 4324
rect 6932 3738 6960 6258
rect 8128 6236 8156 9386
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8220 8090 8248 8230
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8312 7410 8340 9982
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8404 9450 8432 9930
rect 8588 9722 8616 10474
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8680 9518 8708 10406
rect 8772 10130 8800 12406
rect 9140 11898 9168 12786
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9600 10674 9628 12854
rect 10060 12434 10088 13246
rect 10796 12918 10824 13262
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 10060 12406 10180 12434
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9876 11898 9904 12242
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9968 11830 9996 12174
rect 10060 11830 10088 12174
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 10060 11694 10088 11766
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9692 11286 9720 11494
rect 9784 11354 9812 11562
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 10060 10810 10088 11630
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 8760 10124 8812 10130
rect 8760 10066 8812 10072
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8404 9042 8432 9386
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8588 7954 8616 8298
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8588 7546 8616 7890
rect 8680 7546 8708 8230
rect 8864 7886 8892 10610
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 9048 7342 9076 8910
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 8208 6248 8260 6254
rect 8128 6208 8208 6236
rect 8208 6190 8260 6196
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7116 5370 7144 5646
rect 8588 5370 8616 5714
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 9232 5098 9260 9522
rect 9324 8022 9352 10134
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9416 9586 9444 10066
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9508 8906 9536 9454
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9600 9178 9628 9318
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9692 9042 9720 9862
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9600 8498 9720 8514
rect 9600 8492 9732 8498
rect 9600 8486 9680 8492
rect 9312 8016 9364 8022
rect 9312 7958 9364 7964
rect 9600 7886 9628 8486
rect 9680 8434 9732 8440
rect 9784 8362 9812 9522
rect 9876 9110 9904 10542
rect 10152 10062 10180 12406
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10704 11150 10732 11630
rect 10796 11286 10824 12854
rect 11072 12850 11100 13126
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10428 10810 10456 10950
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10888 10606 10916 11494
rect 11072 10606 11100 12786
rect 11164 11286 11192 13382
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 10244 10266 10272 10406
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9968 7954 9996 8230
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 10152 7818 10180 9998
rect 11072 9654 11100 10406
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 11072 9042 11100 9590
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9784 7342 9812 7686
rect 10244 7410 10272 8978
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10428 8090 10456 8230
rect 10704 8090 10732 8774
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10796 8022 10824 8230
rect 10784 8016 10836 8022
rect 10784 7958 10836 7964
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10796 7342 10824 7958
rect 10980 7886 11008 8298
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 9416 6458 9444 7278
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9508 5778 9536 6122
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9220 5092 9272 5098
rect 9220 5034 9272 5040
rect 9324 4146 9352 5646
rect 9404 5160 9456 5166
rect 9508 5148 9536 5714
rect 9456 5120 9536 5148
rect 9404 5102 9456 5108
rect 9600 4282 9628 7142
rect 10796 7002 10824 7278
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10600 6928 10652 6934
rect 10600 6870 10652 6876
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 10060 6322 10088 6666
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9784 5914 9812 6054
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 10244 5778 10272 6190
rect 10232 5772 10284 5778
rect 10232 5714 10284 5720
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10244 5216 10272 5714
rect 10324 5228 10376 5234
rect 10244 5188 10324 5216
rect 10324 5170 10376 5176
rect 9588 4276 9640 4282
rect 9588 4218 9640 4224
rect 10336 4146 10364 5170
rect 10428 5166 10456 5714
rect 10612 5370 10640 6870
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10980 6458 11008 6734
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 7024 3602 7052 3878
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6491 3292 6787 3312
rect 6547 3290 6571 3292
rect 6627 3290 6651 3292
rect 6707 3290 6731 3292
rect 6569 3238 6571 3290
rect 6633 3238 6645 3290
rect 6707 3238 6709 3290
rect 6547 3236 6571 3238
rect 6627 3236 6651 3238
rect 6707 3236 6731 3238
rect 6491 3216 6787 3236
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 11256 2582 11284 14758
rect 11532 14482 11560 16594
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 11624 14414 11652 17546
rect 11716 17202 11744 18702
rect 11808 17542 11836 19246
rect 12026 19068 12322 19088
rect 12082 19066 12106 19068
rect 12162 19066 12186 19068
rect 12242 19066 12266 19068
rect 12104 19014 12106 19066
rect 12168 19014 12180 19066
rect 12242 19014 12244 19066
rect 12082 19012 12106 19014
rect 12162 19012 12186 19014
rect 12242 19012 12266 19014
rect 12026 18992 12322 19012
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12254 18592 12310 18601
rect 12254 18527 12310 18536
rect 12268 18358 12296 18527
rect 12452 18426 12480 18702
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12360 18204 12388 18362
rect 12440 18216 12492 18222
rect 12360 18176 12440 18204
rect 12440 18158 12492 18164
rect 12026 17980 12322 18000
rect 12082 17978 12106 17980
rect 12162 17978 12186 17980
rect 12242 17978 12266 17980
rect 12104 17926 12106 17978
rect 12168 17926 12180 17978
rect 12242 17926 12244 17978
rect 12082 17924 12106 17926
rect 12162 17924 12186 17926
rect 12242 17924 12266 17926
rect 12026 17904 12322 17924
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11900 16794 11928 17682
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12026 16892 12322 16912
rect 12082 16890 12106 16892
rect 12162 16890 12186 16892
rect 12242 16890 12266 16892
rect 12104 16838 12106 16890
rect 12168 16838 12180 16890
rect 12242 16838 12244 16890
rect 12082 16836 12106 16838
rect 12162 16836 12186 16838
rect 12242 16836 12266 16838
rect 12026 16816 12322 16836
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11624 13954 11652 14350
rect 11532 13926 11652 13954
rect 11532 13190 11560 13926
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11624 13394 11652 13806
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11348 9722 11376 10066
rect 11532 10062 11560 10542
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11336 9716 11388 9722
rect 11336 9658 11388 9664
rect 11440 9450 11468 9998
rect 11428 9444 11480 9450
rect 11428 9386 11480 9392
rect 11336 8560 11388 8566
rect 11336 8502 11388 8508
rect 11348 6866 11376 8502
rect 11532 8498 11560 9998
rect 11624 9042 11652 13330
rect 11808 11558 11836 15302
rect 11900 14958 11928 16730
rect 12360 16658 12388 17478
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12440 17060 12492 17066
rect 12440 17002 12492 17008
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12452 15910 12480 17002
rect 12544 16794 12572 17070
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12026 15804 12322 15824
rect 12082 15802 12106 15804
rect 12162 15802 12186 15804
rect 12242 15802 12266 15804
rect 12104 15750 12106 15802
rect 12168 15750 12180 15802
rect 12242 15750 12244 15802
rect 12082 15748 12106 15750
rect 12162 15748 12186 15750
rect 12242 15748 12266 15750
rect 12026 15728 12322 15748
rect 12636 15314 12664 22066
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 12808 21344 12860 21350
rect 12808 21286 12860 21292
rect 12820 21078 12848 21286
rect 12808 21072 12860 21078
rect 12808 21014 12860 21020
rect 12820 19922 12848 21014
rect 12912 20806 12940 21422
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 12912 19786 12940 20742
rect 13188 20398 13216 22578
rect 13360 22568 13412 22574
rect 13360 22510 13412 22516
rect 13372 22098 13400 22510
rect 13360 22092 13412 22098
rect 13360 22034 13412 22040
rect 13452 20528 13504 20534
rect 13452 20470 13504 20476
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 13176 20392 13228 20398
rect 13176 20334 13228 20340
rect 12992 20256 13044 20262
rect 12992 20198 13044 20204
rect 12900 19780 12952 19786
rect 12900 19722 12952 19728
rect 12912 19378 12940 19722
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 12728 18290 12756 18702
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12820 18222 12848 18566
rect 12900 18420 12952 18426
rect 12900 18362 12952 18368
rect 12808 18216 12860 18222
rect 12808 18158 12860 18164
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12728 17678 12756 18022
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12728 15366 12756 16594
rect 12820 15434 12848 16934
rect 12912 16182 12940 18362
rect 13004 17746 13032 20198
rect 13188 19514 13216 20334
rect 13268 20324 13320 20330
rect 13268 20266 13320 20272
rect 13176 19508 13228 19514
rect 13176 19450 13228 19456
rect 13280 19334 13308 20266
rect 13188 19306 13308 19334
rect 13464 19310 13492 20470
rect 13556 19514 13584 20470
rect 13648 20398 13676 23462
rect 13832 22642 13860 23582
rect 14200 23322 14228 26930
rect 14292 26840 14320 35022
rect 14372 31952 14424 31958
rect 14372 31894 14424 31900
rect 14384 31142 14412 31894
rect 14372 31136 14424 31142
rect 14372 31078 14424 31084
rect 14384 30802 14412 31078
rect 14372 30796 14424 30802
rect 14372 30738 14424 30744
rect 14384 29714 14412 30738
rect 14372 29708 14424 29714
rect 14372 29650 14424 29656
rect 14476 26908 14504 35090
rect 15292 34944 15344 34950
rect 15292 34886 15344 34892
rect 14740 33380 14792 33386
rect 14740 33322 14792 33328
rect 14752 31754 14780 33322
rect 14832 32972 14884 32978
rect 14832 32914 14884 32920
rect 14844 32570 14872 32914
rect 15200 32904 15252 32910
rect 15200 32846 15252 32852
rect 14832 32564 14884 32570
rect 14832 32506 14884 32512
rect 15212 32366 15240 32846
rect 15304 32434 15332 34886
rect 15476 33312 15528 33318
rect 15476 33254 15528 33260
rect 15292 32428 15344 32434
rect 15292 32370 15344 32376
rect 15200 32360 15252 32366
rect 15200 32302 15252 32308
rect 15212 32026 15240 32302
rect 15200 32020 15252 32026
rect 15200 31962 15252 31968
rect 15108 31884 15160 31890
rect 15108 31826 15160 31832
rect 14752 31726 14872 31754
rect 14556 28960 14608 28966
rect 14556 28902 14608 28908
rect 14648 28960 14700 28966
rect 14648 28902 14700 28908
rect 14568 28762 14596 28902
rect 14660 28762 14688 28902
rect 14556 28756 14608 28762
rect 14556 28698 14608 28704
rect 14648 28756 14700 28762
rect 14648 28698 14700 28704
rect 14556 27872 14608 27878
rect 14556 27814 14608 27820
rect 14568 27674 14596 27814
rect 14556 27668 14608 27674
rect 14556 27610 14608 27616
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 14476 26880 14688 26908
rect 14292 26812 14504 26840
rect 14372 24676 14424 24682
rect 14372 24618 14424 24624
rect 14188 23316 14240 23322
rect 14188 23258 14240 23264
rect 14384 23118 14412 24618
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 14372 22500 14424 22506
rect 14372 22442 14424 22448
rect 13820 22160 13872 22166
rect 13820 22102 13872 22108
rect 13832 21486 13860 22102
rect 14384 21554 14412 22442
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 14004 21412 14056 21418
rect 14004 21354 14056 21360
rect 14016 20398 14044 21354
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 14004 20392 14056 20398
rect 14004 20334 14056 20340
rect 13544 19508 13596 19514
rect 13544 19450 13596 19456
rect 12992 17740 13044 17746
rect 12992 17682 13044 17688
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 13096 17134 13124 17478
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 12900 16176 12952 16182
rect 12900 16118 12952 16124
rect 13188 15910 13216 19306
rect 13360 19304 13412 19310
rect 13358 19272 13360 19281
rect 13452 19304 13504 19310
rect 13412 19272 13414 19281
rect 13452 19246 13504 19252
rect 13358 19207 13414 19216
rect 13372 18834 13400 19207
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 13280 16658 13308 18158
rect 13464 17082 13492 19246
rect 13556 18766 13584 19450
rect 13648 19378 13676 20334
rect 13912 20256 13964 20262
rect 13912 20198 13964 20204
rect 13820 19440 13872 19446
rect 13820 19382 13872 19388
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 13636 18828 13688 18834
rect 13688 18788 13768 18816
rect 13636 18770 13688 18776
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 13740 18222 13768 18788
rect 13728 18216 13780 18222
rect 13728 18158 13780 18164
rect 13740 17678 13768 18158
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 13648 17134 13676 17478
rect 13740 17270 13768 17614
rect 13728 17264 13780 17270
rect 13728 17206 13780 17212
rect 13636 17128 13688 17134
rect 13464 17066 13584 17082
rect 13636 17070 13688 17076
rect 13464 17060 13596 17066
rect 13464 17054 13544 17060
rect 13544 17002 13596 17008
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13464 16658 13492 16934
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13556 16522 13584 17002
rect 13544 16516 13596 16522
rect 13544 16458 13596 16464
rect 13648 16114 13676 17070
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 12912 15570 12940 15846
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12452 15286 12664 15314
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 12026 14716 12322 14736
rect 12082 14714 12106 14716
rect 12162 14714 12186 14716
rect 12242 14714 12266 14716
rect 12104 14662 12106 14714
rect 12168 14662 12180 14714
rect 12242 14662 12244 14714
rect 12082 14660 12106 14662
rect 12162 14660 12186 14662
rect 12242 14660 12266 14662
rect 12026 14640 12322 14660
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12268 13870 12296 14418
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 12026 13628 12322 13648
rect 12082 13626 12106 13628
rect 12162 13626 12186 13628
rect 12242 13626 12266 13628
rect 12104 13574 12106 13626
rect 12168 13574 12180 13626
rect 12242 13574 12244 13626
rect 12082 13572 12106 13574
rect 12162 13572 12186 13574
rect 12242 13572 12266 13574
rect 12026 13552 12322 13572
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12026 12540 12322 12560
rect 12082 12538 12106 12540
rect 12162 12538 12186 12540
rect 12242 12538 12266 12540
rect 12104 12486 12106 12538
rect 12168 12486 12180 12538
rect 12242 12486 12244 12538
rect 12082 12484 12106 12486
rect 12162 12484 12186 12486
rect 12242 12484 12266 12486
rect 12026 12464 12322 12484
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 12026 11452 12322 11472
rect 12082 11450 12106 11452
rect 12162 11450 12186 11452
rect 12242 11450 12266 11452
rect 12104 11398 12106 11450
rect 12168 11398 12180 11450
rect 12242 11398 12244 11450
rect 12082 11396 12106 11398
rect 12162 11396 12186 11398
rect 12242 11396 12266 11398
rect 12026 11376 12322 11396
rect 12360 10810 12388 12718
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11900 9926 11928 10542
rect 12026 10364 12322 10384
rect 12082 10362 12106 10364
rect 12162 10362 12186 10364
rect 12242 10362 12266 10364
rect 12104 10310 12106 10362
rect 12168 10310 12180 10362
rect 12242 10310 12244 10362
rect 12082 10308 12106 10310
rect 12162 10308 12186 10310
rect 12242 10308 12266 10310
rect 12026 10288 12322 10308
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11624 6798 11652 8978
rect 11900 8430 11928 9862
rect 12026 9276 12322 9296
rect 12082 9274 12106 9276
rect 12162 9274 12186 9276
rect 12242 9274 12266 9276
rect 12104 9222 12106 9274
rect 12168 9222 12180 9274
rect 12242 9222 12244 9274
rect 12082 9220 12106 9222
rect 12162 9220 12186 9222
rect 12242 9220 12266 9222
rect 12026 9200 12322 9220
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 12026 8188 12322 8208
rect 12082 8186 12106 8188
rect 12162 8186 12186 8188
rect 12242 8186 12266 8188
rect 12104 8134 12106 8186
rect 12168 8134 12180 8186
rect 12242 8134 12244 8186
rect 12082 8132 12106 8134
rect 12162 8132 12186 8134
rect 12242 8132 12266 8134
rect 12026 8112 12322 8132
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11992 7342 12020 7686
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11808 5846 11836 7142
rect 12026 7100 12322 7120
rect 12082 7098 12106 7100
rect 12162 7098 12186 7100
rect 12242 7098 12266 7100
rect 12104 7046 12106 7098
rect 12168 7046 12180 7098
rect 12242 7046 12244 7098
rect 12082 7044 12106 7046
rect 12162 7044 12186 7046
rect 12242 7044 12266 7046
rect 12026 7024 12322 7044
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12026 6012 12322 6032
rect 12082 6010 12106 6012
rect 12162 6010 12186 6012
rect 12242 6010 12266 6012
rect 12104 5958 12106 6010
rect 12168 5958 12180 6010
rect 12242 5958 12244 6010
rect 12082 5956 12106 5958
rect 12162 5956 12186 5958
rect 12242 5956 12266 5958
rect 12026 5936 12322 5956
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 12360 5710 12388 6598
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12026 4924 12322 4944
rect 12082 4922 12106 4924
rect 12162 4922 12186 4924
rect 12242 4922 12266 4924
rect 12104 4870 12106 4922
rect 12168 4870 12180 4922
rect 12242 4870 12244 4922
rect 12082 4868 12106 4870
rect 12162 4868 12186 4870
rect 12242 4868 12266 4870
rect 12026 4848 12322 4868
rect 12026 3836 12322 3856
rect 12082 3834 12106 3836
rect 12162 3834 12186 3836
rect 12242 3834 12266 3836
rect 12104 3782 12106 3834
rect 12168 3782 12180 3834
rect 12242 3782 12244 3834
rect 12082 3780 12106 3782
rect 12162 3780 12186 3782
rect 12242 3780 12266 3782
rect 12026 3760 12322 3780
rect 12026 2748 12322 2768
rect 12082 2746 12106 2748
rect 12162 2746 12186 2748
rect 12242 2746 12266 2748
rect 12104 2694 12106 2746
rect 12168 2694 12180 2746
rect 12242 2694 12244 2746
rect 12082 2692 12106 2694
rect 12162 2692 12186 2694
rect 12242 2692 12266 2694
rect 12026 2672 12322 2692
rect 12452 2650 12480 15286
rect 12820 14634 12848 15370
rect 13096 14958 13124 15574
rect 13372 15570 13400 15982
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 12728 14618 13032 14634
rect 12716 14612 13032 14618
rect 12768 14606 13032 14612
rect 12716 14554 12768 14560
rect 12808 14544 12860 14550
rect 12808 14486 12860 14492
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12636 12986 12664 14418
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12728 13530 12756 14214
rect 12820 13920 12848 14486
rect 12900 13932 12952 13938
rect 12820 13892 12900 13920
rect 12820 13530 12848 13892
rect 12900 13874 12952 13880
rect 13004 13870 13032 14606
rect 13096 14414 13124 14894
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 12992 13864 13044 13870
rect 12992 13806 13044 13812
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12820 12782 12848 13466
rect 12912 13326 12940 13670
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12820 11898 12848 12718
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12808 10192 12860 10198
rect 12808 10134 12860 10140
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12544 9178 12572 9318
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12820 9042 12848 10134
rect 12912 9586 12940 12786
rect 13096 12306 13124 13126
rect 13188 12850 13216 14010
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 13096 11558 13124 12242
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 13280 11354 13308 12038
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 13280 10606 13308 11018
rect 13372 10810 13400 15506
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13464 14958 13492 15438
rect 13648 15026 13676 16050
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13740 15570 13768 15846
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13636 15020 13688 15026
rect 13636 14962 13688 14968
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13464 14550 13492 14894
rect 13452 14544 13504 14550
rect 13452 14486 13504 14492
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13556 13870 13584 14214
rect 13648 14074 13676 14962
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13556 13462 13584 13806
rect 13544 13456 13596 13462
rect 13544 13398 13596 13404
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13648 12918 13676 13330
rect 13636 12912 13688 12918
rect 13636 12854 13688 12860
rect 13832 12850 13860 19382
rect 13924 19310 13952 20198
rect 14016 19394 14044 20334
rect 14096 20256 14148 20262
rect 14096 20198 14148 20204
rect 14108 19922 14136 20198
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 14016 19366 14136 19394
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 14004 19236 14056 19242
rect 14004 19178 14056 19184
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 13924 16658 13952 18770
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13924 15910 13952 16594
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13924 12782 13952 13670
rect 14016 12986 14044 19178
rect 14108 16250 14136 19366
rect 14096 16244 14148 16250
rect 14096 16186 14148 16192
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13464 11218 13492 12242
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13360 10804 13412 10810
rect 13360 10746 13412 10752
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12636 7954 12664 8230
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12728 6866 12756 7210
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12820 6390 12848 8978
rect 12912 8362 12940 9522
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12912 7954 12940 8298
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 13004 8090 13032 8230
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 13188 6866 13216 10474
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13280 10266 13308 10406
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13280 9042 13308 10202
rect 13464 10130 13492 11154
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13280 6934 13308 7278
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 13188 6458 13216 6802
rect 13372 6730 13400 9522
rect 13464 9518 13492 10066
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 13464 9178 13492 9454
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13464 8090 13492 8230
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13464 7410 13492 8026
rect 13556 7970 13584 10610
rect 13648 9586 13676 11698
rect 14372 11620 14424 11626
rect 14372 11562 14424 11568
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13740 11218 13768 11494
rect 14096 11280 14148 11286
rect 14096 11222 14148 11228
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13740 10606 13768 11154
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 14108 10538 14136 11222
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 14200 10606 14228 11018
rect 14384 10810 14412 11562
rect 14476 11558 14504 26812
rect 14556 26444 14608 26450
rect 14556 26386 14608 26392
rect 14568 26042 14596 26386
rect 14556 26036 14608 26042
rect 14556 25978 14608 25984
rect 14556 25764 14608 25770
rect 14556 25706 14608 25712
rect 14568 24206 14596 25706
rect 14556 24200 14608 24206
rect 14556 24142 14608 24148
rect 14568 23662 14596 24142
rect 14556 23656 14608 23662
rect 14556 23598 14608 23604
rect 14556 21004 14608 21010
rect 14556 20946 14608 20952
rect 14568 16658 14596 20946
rect 14660 20618 14688 26880
rect 14752 26518 14780 27406
rect 14740 26512 14792 26518
rect 14740 26454 14792 26460
rect 14740 23316 14792 23322
rect 14740 23258 14792 23264
rect 14752 21554 14780 23258
rect 14844 21894 14872 31726
rect 15120 31482 15148 31826
rect 15108 31476 15160 31482
rect 15108 31418 15160 31424
rect 15292 31204 15344 31210
rect 15292 31146 15344 31152
rect 14924 30932 14976 30938
rect 14924 30874 14976 30880
rect 14936 30190 14964 30874
rect 15304 30326 15332 31146
rect 15292 30320 15344 30326
rect 15292 30262 15344 30268
rect 14924 30184 14976 30190
rect 14924 30126 14976 30132
rect 15016 28960 15068 28966
rect 15016 28902 15068 28908
rect 15028 28014 15056 28902
rect 15016 28008 15068 28014
rect 15016 27950 15068 27956
rect 15028 27674 15056 27950
rect 15016 27668 15068 27674
rect 15016 27610 15068 27616
rect 15016 27532 15068 27538
rect 15016 27474 15068 27480
rect 14924 26920 14976 26926
rect 14924 26862 14976 26868
rect 14936 25294 14964 26862
rect 15028 26042 15056 27474
rect 15108 27396 15160 27402
rect 15108 27338 15160 27344
rect 15016 26036 15068 26042
rect 15016 25978 15068 25984
rect 14924 25288 14976 25294
rect 14924 25230 14976 25236
rect 15028 24954 15056 25978
rect 15016 24948 15068 24954
rect 15016 24890 15068 24896
rect 14924 24880 14976 24886
rect 14924 24822 14976 24828
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14740 21548 14792 21554
rect 14740 21490 14792 21496
rect 14936 20942 14964 24822
rect 15016 23180 15068 23186
rect 15016 23122 15068 23128
rect 15028 22778 15056 23122
rect 15016 22772 15068 22778
rect 15016 22714 15068 22720
rect 15016 21480 15068 21486
rect 15016 21422 15068 21428
rect 15028 21146 15056 21422
rect 15016 21140 15068 21146
rect 15016 21082 15068 21088
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 14660 20590 14780 20618
rect 14648 19440 14700 19446
rect 14648 19382 14700 19388
rect 14660 19281 14688 19382
rect 14646 19272 14702 19281
rect 14646 19207 14702 19216
rect 14660 17746 14688 19207
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 14660 16250 14688 17682
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14476 11218 14504 11494
rect 14464 11212 14516 11218
rect 14464 11154 14516 11160
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14096 10532 14148 10538
rect 14096 10474 14148 10480
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13648 9178 13676 9318
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13556 7942 13676 7970
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13360 6724 13412 6730
rect 13360 6666 13412 6672
rect 13464 6458 13492 7346
rect 13556 7002 13584 7822
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13648 6866 13676 7942
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13832 6882 13860 7278
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13740 6854 13860 6882
rect 13544 6724 13596 6730
rect 13544 6666 13596 6672
rect 13556 6458 13584 6666
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 12808 6384 12860 6390
rect 12808 6326 12860 6332
rect 13648 6322 13676 6802
rect 13740 6390 13768 6854
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12636 5914 12664 6190
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 13096 5846 13124 6122
rect 13084 5840 13136 5846
rect 13084 5782 13136 5788
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13372 5166 13400 5510
rect 13648 5370 13676 6258
rect 14016 6254 14044 7142
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 13740 4826 13768 5782
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13004 4146 13032 4762
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13740 4010 13768 4762
rect 14660 4282 14688 12582
rect 14752 10266 14780 20590
rect 14832 20256 14884 20262
rect 14832 20198 14884 20204
rect 14844 19718 14872 20198
rect 15028 19922 15056 21082
rect 15120 21010 15148 27338
rect 15200 25832 15252 25838
rect 15200 25774 15252 25780
rect 15212 24682 15240 25774
rect 15488 25770 15516 33254
rect 15568 26444 15620 26450
rect 15568 26386 15620 26392
rect 15476 25764 15528 25770
rect 15476 25706 15528 25712
rect 15292 24744 15344 24750
rect 15292 24686 15344 24692
rect 15200 24676 15252 24682
rect 15200 24618 15252 24624
rect 15304 24138 15332 24686
rect 15292 24132 15344 24138
rect 15292 24074 15344 24080
rect 15476 23656 15528 23662
rect 15476 23598 15528 23604
rect 15488 22574 15516 23598
rect 15580 22778 15608 26386
rect 15568 22772 15620 22778
rect 15568 22714 15620 22720
rect 15476 22568 15528 22574
rect 15476 22510 15528 22516
rect 15292 22092 15344 22098
rect 15856 22094 15884 35430
rect 16132 35154 16160 36853
rect 18892 35154 18920 36853
rect 21652 35290 21680 36853
rect 23097 35388 23393 35408
rect 23153 35386 23177 35388
rect 23233 35386 23257 35388
rect 23313 35386 23337 35388
rect 23175 35334 23177 35386
rect 23239 35334 23251 35386
rect 23313 35334 23315 35386
rect 23153 35332 23177 35334
rect 23233 35332 23257 35334
rect 23313 35332 23337 35334
rect 23097 35312 23393 35332
rect 24412 35290 24440 36853
rect 21640 35284 21692 35290
rect 21640 35226 21692 35232
rect 24400 35284 24452 35290
rect 24400 35226 24452 35232
rect 27172 35222 27200 36853
rect 27068 35216 27120 35222
rect 27068 35158 27120 35164
rect 27160 35216 27212 35222
rect 27160 35158 27212 35164
rect 16120 35148 16172 35154
rect 16120 35090 16172 35096
rect 18880 35148 18932 35154
rect 18880 35090 18932 35096
rect 21824 35148 21876 35154
rect 21824 35090 21876 35096
rect 20076 35080 20128 35086
rect 20076 35022 20128 35028
rect 18880 34944 18932 34950
rect 18880 34886 18932 34892
rect 17562 34844 17858 34864
rect 17618 34842 17642 34844
rect 17698 34842 17722 34844
rect 17778 34842 17802 34844
rect 17640 34790 17642 34842
rect 17704 34790 17716 34842
rect 17778 34790 17780 34842
rect 17618 34788 17642 34790
rect 17698 34788 17722 34790
rect 17778 34788 17802 34790
rect 17562 34768 17858 34788
rect 16396 34672 16448 34678
rect 16396 34614 16448 34620
rect 16304 34060 16356 34066
rect 16304 34002 16356 34008
rect 16316 32978 16344 34002
rect 16304 32972 16356 32978
rect 16304 32914 16356 32920
rect 16316 31890 16344 32914
rect 16304 31884 16356 31890
rect 16304 31826 16356 31832
rect 16316 31754 16344 31826
rect 16132 31726 16344 31754
rect 16132 31278 16160 31726
rect 16120 31272 16172 31278
rect 16120 31214 16172 31220
rect 16132 30734 16160 31214
rect 16120 30728 16172 30734
rect 16120 30670 16172 30676
rect 16132 29850 16160 30670
rect 16120 29844 16172 29850
rect 16120 29786 16172 29792
rect 16132 29714 16160 29786
rect 16408 29782 16436 34614
rect 17132 34536 17184 34542
rect 17132 34478 17184 34484
rect 17144 34066 17172 34478
rect 17132 34060 17184 34066
rect 17132 34002 17184 34008
rect 18052 33992 18104 33998
rect 18052 33934 18104 33940
rect 17960 33856 18012 33862
rect 17960 33798 18012 33804
rect 17562 33756 17858 33776
rect 17618 33754 17642 33756
rect 17698 33754 17722 33756
rect 17778 33754 17802 33756
rect 17640 33702 17642 33754
rect 17704 33702 17716 33754
rect 17778 33702 17780 33754
rect 17618 33700 17642 33702
rect 17698 33700 17722 33702
rect 17778 33700 17802 33702
rect 17562 33680 17858 33700
rect 17972 33130 18000 33798
rect 18064 33658 18092 33934
rect 18052 33652 18104 33658
rect 18052 33594 18104 33600
rect 18604 33448 18656 33454
rect 18604 33390 18656 33396
rect 18512 33312 18564 33318
rect 18512 33254 18564 33260
rect 17408 33108 17460 33114
rect 17408 33050 17460 33056
rect 17788 33102 18000 33130
rect 17420 31958 17448 33050
rect 17788 33046 17816 33102
rect 18524 33046 18552 33254
rect 17776 33040 17828 33046
rect 17776 32982 17828 32988
rect 18512 33040 18564 33046
rect 18512 32982 18564 32988
rect 17960 32904 18012 32910
rect 17960 32846 18012 32852
rect 17562 32668 17858 32688
rect 17618 32666 17642 32668
rect 17698 32666 17722 32668
rect 17778 32666 17802 32668
rect 17640 32614 17642 32666
rect 17704 32614 17716 32666
rect 17778 32614 17780 32666
rect 17618 32612 17642 32614
rect 17698 32612 17722 32614
rect 17778 32612 17802 32614
rect 17562 32592 17858 32612
rect 17972 32502 18000 32846
rect 17960 32496 18012 32502
rect 17960 32438 18012 32444
rect 18144 32428 18196 32434
rect 18144 32370 18196 32376
rect 17960 32224 18012 32230
rect 17960 32166 18012 32172
rect 17408 31952 17460 31958
rect 17408 31894 17460 31900
rect 16580 31816 16632 31822
rect 16580 31758 16632 31764
rect 16592 31482 16620 31758
rect 16580 31476 16632 31482
rect 16580 31418 16632 31424
rect 17420 30870 17448 31894
rect 17972 31686 18000 32166
rect 17960 31680 18012 31686
rect 17960 31622 18012 31628
rect 17562 31580 17858 31600
rect 17618 31578 17642 31580
rect 17698 31578 17722 31580
rect 17778 31578 17802 31580
rect 17640 31526 17642 31578
rect 17704 31526 17716 31578
rect 17778 31526 17780 31578
rect 17618 31524 17642 31526
rect 17698 31524 17722 31526
rect 17778 31524 17802 31526
rect 17562 31504 17858 31524
rect 17972 31278 18000 31622
rect 18156 31346 18184 32370
rect 18524 32298 18552 32982
rect 18616 32434 18644 33390
rect 18604 32428 18656 32434
rect 18604 32370 18656 32376
rect 18512 32292 18564 32298
rect 18512 32234 18564 32240
rect 18144 31340 18196 31346
rect 18144 31282 18196 31288
rect 18604 31340 18656 31346
rect 18604 31282 18656 31288
rect 17960 31272 18012 31278
rect 17960 31214 18012 31220
rect 17960 31136 18012 31142
rect 17960 31078 18012 31084
rect 17972 30938 18000 31078
rect 17960 30932 18012 30938
rect 17960 30874 18012 30880
rect 17408 30864 17460 30870
rect 17408 30806 17460 30812
rect 17408 30728 17460 30734
rect 17408 30670 17460 30676
rect 17420 30326 17448 30670
rect 17562 30492 17858 30512
rect 17618 30490 17642 30492
rect 17698 30490 17722 30492
rect 17778 30490 17802 30492
rect 17640 30438 17642 30490
rect 17704 30438 17716 30490
rect 17778 30438 17780 30490
rect 17618 30436 17642 30438
rect 17698 30436 17722 30438
rect 17778 30436 17802 30438
rect 17562 30416 17858 30436
rect 17408 30320 17460 30326
rect 17408 30262 17460 30268
rect 17972 30258 18000 30874
rect 17960 30252 18012 30258
rect 17960 30194 18012 30200
rect 18616 30190 18644 31282
rect 18604 30184 18656 30190
rect 18604 30126 18656 30132
rect 16396 29776 16448 29782
rect 16396 29718 16448 29724
rect 16764 29776 16816 29782
rect 16764 29718 16816 29724
rect 16120 29708 16172 29714
rect 16120 29650 16172 29656
rect 16672 29504 16724 29510
rect 16672 29446 16724 29452
rect 16684 29170 16712 29446
rect 16672 29164 16724 29170
rect 16672 29106 16724 29112
rect 16684 28558 16712 29106
rect 16776 29102 16804 29718
rect 18420 29708 18472 29714
rect 18420 29650 18472 29656
rect 17224 29640 17276 29646
rect 17224 29582 17276 29588
rect 18328 29640 18380 29646
rect 18328 29582 18380 29588
rect 16764 29096 16816 29102
rect 16764 29038 16816 29044
rect 16776 28626 16804 29038
rect 16764 28620 16816 28626
rect 16764 28562 16816 28568
rect 16672 28552 16724 28558
rect 16672 28494 16724 28500
rect 16684 27452 16712 28494
rect 16948 28416 17000 28422
rect 16948 28358 17000 28364
rect 16960 28082 16988 28358
rect 16948 28076 17000 28082
rect 16948 28018 17000 28024
rect 17236 27538 17264 29582
rect 17562 29404 17858 29424
rect 17618 29402 17642 29404
rect 17698 29402 17722 29404
rect 17778 29402 17802 29404
rect 17640 29350 17642 29402
rect 17704 29350 17716 29402
rect 17778 29350 17780 29402
rect 17618 29348 17642 29350
rect 17698 29348 17722 29350
rect 17778 29348 17802 29350
rect 17562 29328 17858 29348
rect 18340 29306 18368 29582
rect 18328 29300 18380 29306
rect 18328 29242 18380 29248
rect 17408 29028 17460 29034
rect 17408 28970 17460 28976
rect 17316 28144 17368 28150
rect 17316 28086 17368 28092
rect 17224 27532 17276 27538
rect 17224 27474 17276 27480
rect 16592 27424 16712 27452
rect 16592 26926 16620 27424
rect 16672 26988 16724 26994
rect 16672 26930 16724 26936
rect 16580 26920 16632 26926
rect 16580 26862 16632 26868
rect 16592 26586 16620 26862
rect 16580 26580 16632 26586
rect 16580 26522 16632 26528
rect 16684 26518 16712 26930
rect 17328 26926 17356 28086
rect 17420 27878 17448 28970
rect 17562 28316 17858 28336
rect 17618 28314 17642 28316
rect 17698 28314 17722 28316
rect 17778 28314 17802 28316
rect 17640 28262 17642 28314
rect 17704 28262 17716 28314
rect 17778 28262 17780 28314
rect 17618 28260 17642 28262
rect 17698 28260 17722 28262
rect 17778 28260 17802 28262
rect 17562 28240 17858 28260
rect 17960 27940 18012 27946
rect 17960 27882 18012 27888
rect 17408 27872 17460 27878
rect 17408 27814 17460 27820
rect 17562 27228 17858 27248
rect 17618 27226 17642 27228
rect 17698 27226 17722 27228
rect 17778 27226 17802 27228
rect 17640 27174 17642 27226
rect 17704 27174 17716 27226
rect 17778 27174 17780 27226
rect 17618 27172 17642 27174
rect 17698 27172 17722 27174
rect 17778 27172 17802 27174
rect 17562 27152 17858 27172
rect 17972 26994 18000 27882
rect 18432 27606 18460 29650
rect 18616 29646 18644 30126
rect 18604 29640 18656 29646
rect 18604 29582 18656 29588
rect 18616 29170 18644 29582
rect 18604 29164 18656 29170
rect 18604 29106 18656 29112
rect 18512 27872 18564 27878
rect 18512 27814 18564 27820
rect 18420 27600 18472 27606
rect 18420 27542 18472 27548
rect 18524 27470 18552 27814
rect 18512 27464 18564 27470
rect 18512 27406 18564 27412
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 17316 26920 17368 26926
rect 17316 26862 17368 26868
rect 18604 26920 18656 26926
rect 18604 26862 18656 26868
rect 16672 26512 16724 26518
rect 16672 26454 16724 26460
rect 17328 26450 17356 26862
rect 17316 26444 17368 26450
rect 17316 26386 17368 26392
rect 17562 26140 17858 26160
rect 17618 26138 17642 26140
rect 17698 26138 17722 26140
rect 17778 26138 17802 26140
rect 17640 26086 17642 26138
rect 17704 26086 17716 26138
rect 17778 26086 17780 26138
rect 17618 26084 17642 26086
rect 17698 26084 17722 26086
rect 17778 26084 17802 26086
rect 17562 26064 17858 26084
rect 16672 25832 16724 25838
rect 16672 25774 16724 25780
rect 17408 25832 17460 25838
rect 17408 25774 17460 25780
rect 17500 25832 17552 25838
rect 17500 25774 17552 25780
rect 16028 25696 16080 25702
rect 16028 25638 16080 25644
rect 16580 25696 16632 25702
rect 16580 25638 16632 25644
rect 16040 24750 16068 25638
rect 16212 25356 16264 25362
rect 16212 25298 16264 25304
rect 16224 24954 16252 25298
rect 16212 24948 16264 24954
rect 16212 24890 16264 24896
rect 16304 24812 16356 24818
rect 16304 24754 16356 24760
rect 16028 24744 16080 24750
rect 16028 24686 16080 24692
rect 16316 24342 16344 24754
rect 16592 24750 16620 25638
rect 16684 25158 16712 25774
rect 16672 25152 16724 25158
rect 16672 25094 16724 25100
rect 17132 25152 17184 25158
rect 17132 25094 17184 25100
rect 16684 24818 16712 25094
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16580 24744 16632 24750
rect 16580 24686 16632 24692
rect 17144 24682 17172 25094
rect 17420 24750 17448 25774
rect 17512 25226 17540 25774
rect 18144 25356 18196 25362
rect 18144 25298 18196 25304
rect 17500 25220 17552 25226
rect 17500 25162 17552 25168
rect 17562 25052 17858 25072
rect 17618 25050 17642 25052
rect 17698 25050 17722 25052
rect 17778 25050 17802 25052
rect 17640 24998 17642 25050
rect 17704 24998 17716 25050
rect 17778 24998 17780 25050
rect 17618 24996 17642 24998
rect 17698 24996 17722 24998
rect 17778 24996 17802 24998
rect 17562 24976 17858 24996
rect 17408 24744 17460 24750
rect 17408 24686 17460 24692
rect 17132 24676 17184 24682
rect 17132 24618 17184 24624
rect 16304 24336 16356 24342
rect 16304 24278 16356 24284
rect 17144 24274 17172 24618
rect 17224 24608 17276 24614
rect 17224 24550 17276 24556
rect 17132 24268 17184 24274
rect 17132 24210 17184 24216
rect 17236 24206 17264 24550
rect 17224 24200 17276 24206
rect 17224 24142 17276 24148
rect 16120 24132 16172 24138
rect 16120 24074 16172 24080
rect 16132 23254 16160 24074
rect 17420 23322 17448 24686
rect 18156 24410 18184 25298
rect 18144 24404 18196 24410
rect 18144 24346 18196 24352
rect 17960 24064 18012 24070
rect 17960 24006 18012 24012
rect 17562 23964 17858 23984
rect 17618 23962 17642 23964
rect 17698 23962 17722 23964
rect 17778 23962 17802 23964
rect 17640 23910 17642 23962
rect 17704 23910 17716 23962
rect 17778 23910 17780 23962
rect 17618 23908 17642 23910
rect 17698 23908 17722 23910
rect 17778 23908 17802 23910
rect 17562 23888 17858 23908
rect 17972 23322 18000 24006
rect 17408 23316 17460 23322
rect 17408 23258 17460 23264
rect 17960 23316 18012 23322
rect 17960 23258 18012 23264
rect 16120 23248 16172 23254
rect 16120 23190 16172 23196
rect 16304 23248 16356 23254
rect 16304 23190 16356 23196
rect 16672 23248 16724 23254
rect 16672 23190 16724 23196
rect 16316 22642 16344 23190
rect 16304 22636 16356 22642
rect 16304 22578 16356 22584
rect 15856 22066 16252 22094
rect 15292 22034 15344 22040
rect 15108 21004 15160 21010
rect 15108 20946 15160 20952
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15016 19916 15068 19922
rect 15016 19858 15068 19864
rect 14832 19712 14884 19718
rect 14832 19654 14884 19660
rect 14924 19712 14976 19718
rect 14924 19654 14976 19660
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 14844 19174 14872 19450
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14936 18986 14964 19654
rect 15014 19272 15070 19281
rect 15014 19207 15016 19216
rect 15068 19207 15070 19216
rect 15016 19178 15068 19184
rect 14844 18958 14964 18986
rect 14844 18290 14872 18958
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 14844 17542 14872 18226
rect 14936 17814 14964 18770
rect 15028 18426 15056 19178
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 15016 18420 15068 18426
rect 15016 18362 15068 18368
rect 15016 18216 15068 18222
rect 15016 18158 15068 18164
rect 14924 17808 14976 17814
rect 14924 17750 14976 17756
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14936 16946 14964 17750
rect 15028 17134 15056 18158
rect 15120 17202 15148 19110
rect 15212 18766 15240 19994
rect 15304 19242 15332 22034
rect 15844 20324 15896 20330
rect 15844 20266 15896 20272
rect 16120 20324 16172 20330
rect 16120 20266 16172 20272
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 15764 19378 15792 19654
rect 15856 19514 15884 20266
rect 16132 19786 16160 20266
rect 16120 19780 16172 19786
rect 16120 19722 16172 19728
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 15844 19508 15896 19514
rect 15844 19450 15896 19456
rect 16040 19446 16068 19654
rect 16028 19440 16080 19446
rect 16028 19382 16080 19388
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15844 19304 15896 19310
rect 15844 19246 15896 19252
rect 15292 19236 15344 19242
rect 15292 19178 15344 19184
rect 15488 18902 15516 19246
rect 15752 19236 15804 19242
rect 15752 19178 15804 19184
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 15764 18426 15792 19178
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15396 17814 15424 18022
rect 15384 17808 15436 17814
rect 15384 17750 15436 17756
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 14936 16918 15056 16946
rect 15028 16726 15056 16918
rect 15120 16794 15148 17138
rect 15108 16788 15160 16794
rect 15108 16730 15160 16736
rect 15016 16720 15068 16726
rect 15016 16662 15068 16668
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 14844 16114 14872 16594
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 15028 13462 15056 14214
rect 15212 13530 15240 17614
rect 15396 17066 15424 17750
rect 15488 17746 15516 18158
rect 15856 18086 15884 19246
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15948 17814 15976 19110
rect 16040 18834 16068 19382
rect 16132 19310 16160 19722
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 16028 18828 16080 18834
rect 16028 18770 16080 18776
rect 15936 17808 15988 17814
rect 15936 17750 15988 17756
rect 16120 17808 16172 17814
rect 16120 17750 16172 17756
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 16132 17202 16160 17750
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 15384 17060 15436 17066
rect 15384 17002 15436 17008
rect 15752 17060 15804 17066
rect 15752 17002 15804 17008
rect 15476 16516 15528 16522
rect 15476 16458 15528 16464
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 15304 14074 15332 14418
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15396 13870 15424 15642
rect 15488 14958 15516 16458
rect 15764 15978 15792 17002
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15948 16046 15976 16390
rect 15936 16040 15988 16046
rect 15936 15982 15988 15988
rect 15752 15972 15804 15978
rect 15752 15914 15804 15920
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15580 15570 15608 15846
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15660 14884 15712 14890
rect 15660 14826 15712 14832
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15016 13456 15068 13462
rect 15016 13398 15068 13404
rect 15212 11898 15240 13466
rect 15292 13456 15344 13462
rect 15396 13410 15424 13670
rect 15344 13404 15424 13410
rect 15292 13398 15424 13404
rect 15304 13382 15424 13398
rect 15396 13326 15424 13382
rect 15488 13326 15516 14350
rect 15672 14074 15700 14826
rect 15764 14482 15792 15302
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15672 13852 15700 14010
rect 15752 13864 15804 13870
rect 15672 13824 15752 13852
rect 15752 13806 15804 13812
rect 16132 13734 16160 17138
rect 16224 15994 16252 22066
rect 16316 20942 16344 22578
rect 16580 22228 16632 22234
rect 16684 22216 16712 23190
rect 17224 23180 17276 23186
rect 17224 23122 17276 23128
rect 16632 22188 16712 22216
rect 16580 22170 16632 22176
rect 16580 22092 16632 22098
rect 16580 22034 16632 22040
rect 16592 22001 16620 22034
rect 16578 21992 16634 22001
rect 16578 21927 16634 21936
rect 16580 21004 16632 21010
rect 16580 20946 16632 20952
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 16316 20466 16344 20878
rect 16304 20460 16356 20466
rect 16304 20402 16356 20408
rect 16592 20058 16620 20946
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16304 19984 16356 19990
rect 16304 19926 16356 19932
rect 16316 18902 16344 19926
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16592 19242 16620 19654
rect 16580 19236 16632 19242
rect 16580 19178 16632 19184
rect 16304 18896 16356 18902
rect 16304 18838 16356 18844
rect 16684 18601 16712 22188
rect 16764 20324 16816 20330
rect 16764 20266 16816 20272
rect 16776 19922 16804 20266
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 17236 18714 17264 23122
rect 17562 22876 17858 22896
rect 17618 22874 17642 22876
rect 17698 22874 17722 22876
rect 17778 22874 17802 22876
rect 17640 22822 17642 22874
rect 17704 22822 17716 22874
rect 17778 22822 17780 22874
rect 17618 22820 17642 22822
rect 17698 22820 17722 22822
rect 17778 22820 17802 22822
rect 17562 22800 17858 22820
rect 17316 22432 17368 22438
rect 17316 22374 17368 22380
rect 17328 20398 17356 22374
rect 18616 22166 18644 26862
rect 18696 26444 18748 26450
rect 18696 26386 18748 26392
rect 18708 23186 18736 26386
rect 18788 26308 18840 26314
rect 18788 26250 18840 26256
rect 18800 25430 18828 26250
rect 18788 25424 18840 25430
rect 18788 25366 18840 25372
rect 18800 24342 18828 25366
rect 18788 24336 18840 24342
rect 18788 24278 18840 24284
rect 18696 23180 18748 23186
rect 18696 23122 18748 23128
rect 18788 22976 18840 22982
rect 18788 22918 18840 22924
rect 18800 22642 18828 22918
rect 18788 22636 18840 22642
rect 18788 22578 18840 22584
rect 18604 22160 18656 22166
rect 18604 22102 18656 22108
rect 17562 21788 17858 21808
rect 17618 21786 17642 21788
rect 17698 21786 17722 21788
rect 17778 21786 17802 21788
rect 17640 21734 17642 21786
rect 17704 21734 17716 21786
rect 17778 21734 17780 21786
rect 17618 21732 17642 21734
rect 17698 21732 17722 21734
rect 17778 21732 17802 21734
rect 17562 21712 17858 21732
rect 17684 21480 17736 21486
rect 17684 21422 17736 21428
rect 17696 21146 17724 21422
rect 18696 21412 18748 21418
rect 18696 21354 18748 21360
rect 18512 21344 18564 21350
rect 18512 21286 18564 21292
rect 17408 21140 17460 21146
rect 17408 21082 17460 21088
rect 17684 21140 17736 21146
rect 17684 21082 17736 21088
rect 17420 20398 17448 21082
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 17562 20700 17858 20720
rect 17618 20698 17642 20700
rect 17698 20698 17722 20700
rect 17778 20698 17802 20700
rect 17640 20646 17642 20698
rect 17704 20646 17716 20698
rect 17778 20646 17780 20698
rect 17618 20644 17642 20646
rect 17698 20644 17722 20646
rect 17778 20644 17802 20646
rect 17562 20624 17858 20644
rect 18340 20398 18368 20742
rect 17316 20392 17368 20398
rect 17316 20334 17368 20340
rect 17408 20392 17460 20398
rect 17408 20334 17460 20340
rect 18328 20392 18380 20398
rect 18328 20334 18380 20340
rect 18420 20256 18472 20262
rect 18420 20198 18472 20204
rect 17316 19916 17368 19922
rect 17316 19858 17368 19864
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17328 19281 17356 19858
rect 17880 19700 17908 19858
rect 17880 19672 18000 19700
rect 17562 19612 17858 19632
rect 17618 19610 17642 19612
rect 17698 19610 17722 19612
rect 17778 19610 17802 19612
rect 17640 19558 17642 19610
rect 17704 19558 17716 19610
rect 17778 19558 17780 19610
rect 17618 19556 17642 19558
rect 17698 19556 17722 19558
rect 17778 19556 17802 19558
rect 17562 19536 17858 19556
rect 17972 19496 18000 19672
rect 17880 19468 18000 19496
rect 17314 19272 17370 19281
rect 17314 19207 17370 19216
rect 17776 19236 17828 19242
rect 17776 19178 17828 19184
rect 17788 18970 17816 19178
rect 17408 18964 17460 18970
rect 17408 18906 17460 18912
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 16868 18698 17264 18714
rect 16856 18692 17264 18698
rect 16908 18686 17264 18692
rect 16856 18634 16908 18640
rect 17040 18624 17092 18630
rect 16670 18592 16726 18601
rect 17040 18566 17092 18572
rect 16670 18527 16726 18536
rect 16684 18358 16712 18527
rect 16672 18352 16724 18358
rect 16672 18294 16724 18300
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16408 16250 16436 16594
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16960 16182 16988 16390
rect 16948 16176 17000 16182
rect 16948 16118 17000 16124
rect 16224 15966 16344 15994
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16224 14958 16252 15846
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 16224 13870 16252 14894
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16120 13728 16172 13734
rect 16316 13682 16344 15966
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16396 15020 16448 15026
rect 16396 14962 16448 14968
rect 16408 13870 16436 14962
rect 16592 14618 16620 15506
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16684 14890 16712 15438
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16120 13670 16172 13676
rect 16224 13654 16344 13682
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14936 10674 14964 10950
rect 15488 10810 15516 12038
rect 15580 11694 15608 12038
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15764 11354 15792 12174
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 15212 9178 15240 10542
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15488 10198 15516 10406
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15476 10192 15528 10198
rect 15476 10134 15528 10140
rect 15580 9518 15608 10202
rect 15672 9722 15700 10610
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15856 9518 15884 11154
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14752 6322 14780 7822
rect 15396 6730 15424 8366
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15476 7948 15528 7954
rect 15476 7890 15528 7896
rect 15488 7546 15516 7890
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15580 7410 15608 8230
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14752 5710 14780 6258
rect 15396 5710 15424 6666
rect 15764 6662 15792 7278
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15580 6254 15608 6598
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15948 5914 15976 6802
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 14752 4690 14780 5646
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 15028 4758 15056 4966
rect 15016 4752 15068 4758
rect 15016 4694 15068 4700
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14752 4146 14780 4626
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 16040 2582 16068 13262
rect 16224 12782 16252 13654
rect 16776 13462 16804 14418
rect 16856 14340 16908 14346
rect 16856 14282 16908 14288
rect 16764 13456 16816 13462
rect 16764 13398 16816 13404
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16316 12986 16344 13330
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16776 11898 16804 12242
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16132 10130 16160 11698
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16408 10470 16436 10746
rect 16488 10736 16540 10742
rect 16488 10678 16540 10684
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 16132 8430 16160 8978
rect 16224 8634 16252 8978
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 16132 8090 16160 8366
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16224 6458 16252 6802
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16120 6180 16172 6186
rect 16120 6122 16172 6128
rect 16132 5778 16160 6122
rect 16224 5846 16252 6394
rect 16212 5840 16264 5846
rect 16212 5782 16264 5788
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 16132 5030 16160 5714
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16316 4758 16344 5170
rect 16304 4752 16356 4758
rect 16304 4694 16356 4700
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 11244 2576 11296 2582
rect 11244 2518 11296 2524
rect 16028 2576 16080 2582
rect 16028 2518 16080 2524
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 480 2372 532 2378
rect 480 2314 532 2320
rect 492 800 520 2314
rect 2792 800 2820 2450
rect 5552 800 5580 2450
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 11060 2372 11112 2378
rect 11060 2314 11112 2320
rect 6491 2204 6787 2224
rect 6547 2202 6571 2204
rect 6627 2202 6651 2204
rect 6707 2202 6731 2204
rect 6569 2150 6571 2202
rect 6633 2150 6645 2202
rect 6707 2150 6709 2202
rect 6547 2148 6571 2150
rect 6627 2148 6651 2150
rect 6707 2148 6731 2150
rect 6491 2128 6787 2148
rect 8312 800 8340 2314
rect 11072 800 11100 2314
rect 13832 800 13860 2450
rect 16132 2446 16160 3334
rect 16408 2774 16436 10406
rect 16500 10266 16528 10678
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16500 9738 16528 10202
rect 16764 10192 16816 10198
rect 16764 10134 16816 10140
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 16500 9710 16620 9738
rect 16592 7818 16620 9710
rect 16684 9178 16712 10066
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16580 7812 16632 7818
rect 16580 7754 16632 7760
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16684 7342 16712 7686
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16776 6866 16804 10134
rect 16868 9654 16896 14282
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16856 9648 16908 9654
rect 16856 9590 16908 9596
rect 16960 8634 16988 10066
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 17052 8430 17080 18566
rect 17236 17882 17264 18686
rect 17420 18426 17448 18906
rect 17880 18698 17908 19468
rect 18052 18896 18104 18902
rect 18052 18838 18104 18844
rect 17868 18692 17920 18698
rect 17868 18634 17920 18640
rect 17562 18524 17858 18544
rect 17618 18522 17642 18524
rect 17698 18522 17722 18524
rect 17778 18522 17802 18524
rect 17640 18470 17642 18522
rect 17704 18470 17716 18522
rect 17778 18470 17780 18522
rect 17618 18468 17642 18470
rect 17698 18468 17722 18470
rect 17778 18468 17802 18470
rect 17562 18448 17858 18468
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17420 17746 17448 18362
rect 18064 18290 18092 18838
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 17408 17740 17460 17746
rect 17408 17682 17460 17688
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 17236 17066 17264 17478
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 17224 17060 17276 17066
rect 17224 17002 17276 17008
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 17144 16114 17172 16934
rect 17236 16658 17264 17002
rect 17328 16726 17356 17138
rect 17420 16794 17448 17682
rect 17562 17436 17858 17456
rect 17618 17434 17642 17436
rect 17698 17434 17722 17436
rect 17778 17434 17802 17436
rect 17640 17382 17642 17434
rect 17704 17382 17716 17434
rect 17778 17382 17780 17434
rect 17618 17380 17642 17382
rect 17698 17380 17722 17382
rect 17778 17380 17802 17382
rect 17562 17360 17858 17380
rect 17408 16788 17460 16794
rect 17408 16730 17460 16736
rect 17316 16720 17368 16726
rect 17316 16662 17368 16668
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 17132 16108 17184 16114
rect 17132 16050 17184 16056
rect 17144 15586 17172 16050
rect 17328 15978 17356 16526
rect 17562 16348 17858 16368
rect 17618 16346 17642 16348
rect 17698 16346 17722 16348
rect 17778 16346 17802 16348
rect 17640 16294 17642 16346
rect 17704 16294 17716 16346
rect 17778 16294 17780 16346
rect 17618 16292 17642 16294
rect 17698 16292 17722 16294
rect 17778 16292 17802 16294
rect 17562 16272 17858 16292
rect 17316 15972 17368 15978
rect 17316 15914 17368 15920
rect 17328 15638 17356 15914
rect 17316 15632 17368 15638
rect 17144 15570 17264 15586
rect 17316 15574 17368 15580
rect 17144 15564 17276 15570
rect 17144 15558 17224 15564
rect 17224 15506 17276 15512
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17880 15450 17908 15506
rect 17880 15422 18000 15450
rect 17408 15360 17460 15366
rect 17408 15302 17460 15308
rect 17420 15162 17448 15302
rect 17562 15260 17858 15280
rect 17618 15258 17642 15260
rect 17698 15258 17722 15260
rect 17778 15258 17802 15260
rect 17640 15206 17642 15258
rect 17704 15206 17716 15258
rect 17778 15206 17780 15258
rect 17618 15204 17642 15206
rect 17698 15204 17722 15206
rect 17778 15204 17802 15206
rect 17562 15184 17858 15204
rect 17972 15162 18000 15422
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17328 14074 17356 14894
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17420 14006 17448 14758
rect 18432 14550 18460 20198
rect 18420 14544 18472 14550
rect 18420 14486 18472 14492
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17562 14172 17858 14192
rect 17618 14170 17642 14172
rect 17698 14170 17722 14172
rect 17778 14170 17802 14172
rect 17640 14118 17642 14170
rect 17704 14118 17716 14170
rect 17778 14118 17780 14170
rect 17618 14116 17642 14118
rect 17698 14116 17722 14118
rect 17778 14116 17802 14118
rect 17562 14096 17858 14116
rect 17408 14000 17460 14006
rect 17408 13942 17460 13948
rect 17420 13394 17448 13942
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17562 13084 17858 13104
rect 17618 13082 17642 13084
rect 17698 13082 17722 13084
rect 17778 13082 17802 13084
rect 17640 13030 17642 13082
rect 17704 13030 17716 13082
rect 17778 13030 17780 13082
rect 17618 13028 17642 13030
rect 17698 13028 17722 13030
rect 17778 13028 17802 13030
rect 17562 13008 17858 13028
rect 17972 12850 18000 14418
rect 18236 14408 18288 14414
rect 18288 14356 18368 14362
rect 18236 14350 18368 14356
rect 18248 14334 18368 14350
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18248 13870 18276 14214
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 18236 13388 18288 13394
rect 18236 13330 18288 13336
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 17684 12776 17736 12782
rect 17684 12718 17736 12724
rect 18052 12776 18104 12782
rect 18248 12764 18276 13330
rect 18052 12718 18104 12724
rect 18156 12736 18276 12764
rect 17696 12442 17724 12718
rect 17960 12708 18012 12714
rect 17960 12650 18012 12656
rect 17972 12442 18000 12650
rect 17684 12436 17736 12442
rect 17684 12378 17736 12384
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17224 12164 17276 12170
rect 17224 12106 17276 12112
rect 17236 11014 17264 12106
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 17144 8634 17172 9862
rect 17236 9178 17264 10542
rect 17328 10198 17356 12242
rect 17562 11996 17858 12016
rect 17618 11994 17642 11996
rect 17698 11994 17722 11996
rect 17778 11994 17802 11996
rect 17640 11942 17642 11994
rect 17704 11942 17716 11994
rect 17778 11942 17780 11994
rect 17618 11940 17642 11942
rect 17698 11940 17722 11942
rect 17778 11940 17802 11942
rect 17562 11920 17858 11940
rect 17408 11008 17460 11014
rect 17408 10950 17460 10956
rect 17316 10192 17368 10198
rect 17316 10134 17368 10140
rect 17420 10130 17448 10950
rect 17562 10908 17858 10928
rect 17618 10906 17642 10908
rect 17698 10906 17722 10908
rect 17778 10906 17802 10908
rect 17640 10854 17642 10906
rect 17704 10854 17716 10906
rect 17778 10854 17780 10906
rect 17618 10852 17642 10854
rect 17698 10852 17722 10854
rect 17778 10852 17802 10854
rect 17562 10832 17858 10852
rect 17972 10130 18000 12242
rect 18064 11354 18092 12718
rect 18156 12374 18184 12736
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 18144 12368 18196 12374
rect 18144 12310 18196 12316
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 18144 11212 18196 11218
rect 18144 11154 18196 11160
rect 18156 10538 18184 11154
rect 18248 10690 18276 12378
rect 18340 12102 18368 14334
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18432 11234 18460 13330
rect 18524 12782 18552 21286
rect 18708 21010 18736 21354
rect 18696 21004 18748 21010
rect 18696 20946 18748 20952
rect 18708 19786 18736 20946
rect 18696 19780 18748 19786
rect 18696 19722 18748 19728
rect 18604 18148 18656 18154
rect 18604 18090 18656 18096
rect 18616 16998 18644 18090
rect 18604 16992 18656 16998
rect 18604 16934 18656 16940
rect 18616 16658 18644 16934
rect 18604 16652 18656 16658
rect 18604 16594 18656 16600
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 18788 14476 18840 14482
rect 18788 14418 18840 14424
rect 18708 13394 18736 14418
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18800 12918 18828 14418
rect 18788 12912 18840 12918
rect 18788 12854 18840 12860
rect 18512 12776 18564 12782
rect 18512 12718 18564 12724
rect 18892 12374 18920 34886
rect 19892 34604 19944 34610
rect 19892 34546 19944 34552
rect 19432 34536 19484 34542
rect 19432 34478 19484 34484
rect 19340 33856 19392 33862
rect 19340 33798 19392 33804
rect 19352 33318 19380 33798
rect 19444 33658 19472 34478
rect 19432 33652 19484 33658
rect 19432 33594 19484 33600
rect 19904 33522 19932 34546
rect 19892 33516 19944 33522
rect 19892 33458 19944 33464
rect 19340 33312 19392 33318
rect 19340 33254 19392 33260
rect 19800 33312 19852 33318
rect 19800 33254 19852 33260
rect 19812 32910 19840 33254
rect 19800 32904 19852 32910
rect 19800 32846 19852 32852
rect 19156 32836 19208 32842
rect 19156 32778 19208 32784
rect 19168 32366 19196 32778
rect 19904 32774 19932 33458
rect 19892 32768 19944 32774
rect 19892 32710 19944 32716
rect 19340 32496 19392 32502
rect 19340 32438 19392 32444
rect 19156 32360 19208 32366
rect 19156 32302 19208 32308
rect 19064 31136 19116 31142
rect 19064 31078 19116 31084
rect 19076 28626 19104 31078
rect 19156 30252 19208 30258
rect 19156 30194 19208 30200
rect 19168 29170 19196 30194
rect 19156 29164 19208 29170
rect 19156 29106 19208 29112
rect 19064 28620 19116 28626
rect 19064 28562 19116 28568
rect 18972 28484 19024 28490
rect 18972 28426 19024 28432
rect 18984 26586 19012 28426
rect 19168 28082 19196 29106
rect 19352 28694 19380 32438
rect 19616 31204 19668 31210
rect 19616 31146 19668 31152
rect 19628 30734 19656 31146
rect 19616 30728 19668 30734
rect 19616 30670 19668 30676
rect 19628 30054 19656 30670
rect 19616 30048 19668 30054
rect 19616 29990 19668 29996
rect 19628 29102 19656 29990
rect 19616 29096 19668 29102
rect 19616 29038 19668 29044
rect 19340 28688 19392 28694
rect 19340 28630 19392 28636
rect 19340 28416 19392 28422
rect 19340 28358 19392 28364
rect 19156 28076 19208 28082
rect 19156 28018 19208 28024
rect 19168 27878 19196 28018
rect 19064 27872 19116 27878
rect 19064 27814 19116 27820
rect 19156 27872 19208 27878
rect 19156 27814 19208 27820
rect 19076 27334 19104 27814
rect 19064 27328 19116 27334
rect 19064 27270 19116 27276
rect 19076 26926 19104 27270
rect 19064 26920 19116 26926
rect 19064 26862 19116 26868
rect 18972 26580 19024 26586
rect 18972 26522 19024 26528
rect 19076 26450 19104 26862
rect 19064 26444 19116 26450
rect 19064 26386 19116 26392
rect 19156 25832 19208 25838
rect 19156 25774 19208 25780
rect 19168 25294 19196 25774
rect 19156 25288 19208 25294
rect 19156 25230 19208 25236
rect 19168 24818 19196 25230
rect 19156 24812 19208 24818
rect 19156 24754 19208 24760
rect 19352 23186 19380 28358
rect 19432 27532 19484 27538
rect 19432 27474 19484 27480
rect 19800 27532 19852 27538
rect 19800 27474 19852 27480
rect 19444 26994 19472 27474
rect 19432 26988 19484 26994
rect 19432 26930 19484 26936
rect 19444 26586 19472 26930
rect 19432 26580 19484 26586
rect 19432 26522 19484 26528
rect 19432 24676 19484 24682
rect 19432 24618 19484 24624
rect 19444 23866 19472 24618
rect 19524 24608 19576 24614
rect 19524 24550 19576 24556
rect 19432 23860 19484 23866
rect 19432 23802 19484 23808
rect 19536 23202 19564 24550
rect 19616 23520 19668 23526
rect 19616 23462 19668 23468
rect 19628 23254 19656 23462
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19444 23174 19564 23202
rect 19616 23248 19668 23254
rect 19616 23190 19668 23196
rect 19444 22658 19472 23174
rect 19524 23112 19576 23118
rect 19524 23054 19576 23060
rect 19536 22778 19564 23054
rect 19524 22772 19576 22778
rect 19524 22714 19576 22720
rect 19628 22710 19656 23190
rect 19352 22630 19472 22658
rect 19616 22704 19668 22710
rect 19616 22646 19668 22652
rect 19352 22506 19380 22630
rect 19432 22568 19484 22574
rect 19432 22510 19484 22516
rect 19340 22500 19392 22506
rect 19340 22442 19392 22448
rect 19444 22030 19472 22510
rect 19708 22500 19760 22506
rect 19708 22442 19760 22448
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19720 21554 19748 22442
rect 19708 21548 19760 21554
rect 19708 21490 19760 21496
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19064 20868 19116 20874
rect 19064 20810 19116 20816
rect 18972 20800 19024 20806
rect 18972 20742 19024 20748
rect 18984 19990 19012 20742
rect 19076 20262 19104 20810
rect 19444 20602 19472 20878
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 19076 20058 19104 20198
rect 19064 20052 19116 20058
rect 19064 19994 19116 20000
rect 18972 19984 19024 19990
rect 18972 19926 19024 19932
rect 19812 19258 19840 27474
rect 19984 22568 20036 22574
rect 19984 22510 20036 22516
rect 19892 22432 19944 22438
rect 19892 22374 19944 22380
rect 19904 19310 19932 22374
rect 19996 21690 20024 22510
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 19536 19230 19840 19258
rect 19892 19304 19944 19310
rect 19892 19246 19944 19252
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 18984 18086 19012 18702
rect 19536 18698 19564 19230
rect 19800 19168 19852 19174
rect 19800 19110 19852 19116
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 19064 18624 19116 18630
rect 19064 18566 19116 18572
rect 19076 18290 19104 18566
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 19628 17542 19656 18702
rect 19720 18358 19748 18770
rect 19812 18766 19840 19110
rect 19904 18970 19932 19246
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19890 18864 19946 18873
rect 19890 18799 19892 18808
rect 19944 18799 19946 18808
rect 19892 18770 19944 18776
rect 19800 18760 19852 18766
rect 19800 18702 19852 18708
rect 19904 18426 19932 18770
rect 19892 18420 19944 18426
rect 19892 18362 19944 18368
rect 19708 18352 19760 18358
rect 19708 18294 19760 18300
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19996 17134 20024 17478
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 18972 17060 19024 17066
rect 18972 17002 19024 17008
rect 18984 16250 19012 17002
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 19524 16244 19576 16250
rect 19524 16186 19576 16192
rect 19536 15978 19564 16186
rect 19812 16114 19840 16934
rect 19996 16454 20024 17070
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 19996 16182 20024 16390
rect 19984 16176 20036 16182
rect 19984 16118 20036 16124
rect 19800 16108 19852 16114
rect 19800 16050 19852 16056
rect 19524 15972 19576 15978
rect 19524 15914 19576 15920
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 19076 14822 19104 15438
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 18972 14476 19024 14482
rect 18972 14418 19024 14424
rect 18984 14006 19012 14418
rect 19076 14346 19104 14758
rect 19984 14476 20036 14482
rect 19984 14418 20036 14424
rect 19064 14340 19116 14346
rect 19064 14282 19116 14288
rect 19996 14074 20024 14418
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 18972 14000 19024 14006
rect 18972 13942 19024 13948
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18880 12368 18932 12374
rect 18880 12310 18932 12316
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18524 11286 18552 11630
rect 18340 11206 18460 11234
rect 18512 11280 18564 11286
rect 18512 11222 18564 11228
rect 18340 10810 18368 11206
rect 18420 11076 18472 11082
rect 18420 11018 18472 11024
rect 18328 10804 18380 10810
rect 18328 10746 18380 10752
rect 18248 10662 18368 10690
rect 18432 10674 18460 11018
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 18144 10532 18196 10538
rect 18144 10474 18196 10480
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17328 9518 17356 9998
rect 17562 9820 17858 9840
rect 17618 9818 17642 9820
rect 17698 9818 17722 9820
rect 17778 9818 17802 9820
rect 17640 9766 17642 9818
rect 17704 9766 17716 9818
rect 17778 9766 17780 9818
rect 17618 9764 17642 9766
rect 17698 9764 17722 9766
rect 17778 9764 17802 9766
rect 17562 9744 17858 9764
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17224 9036 17276 9042
rect 17224 8978 17276 8984
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17040 8424 17092 8430
rect 17040 8366 17092 8372
rect 17236 8362 17264 8978
rect 17562 8732 17858 8752
rect 17618 8730 17642 8732
rect 17698 8730 17722 8732
rect 17778 8730 17802 8732
rect 17640 8678 17642 8730
rect 17704 8678 17716 8730
rect 17778 8678 17780 8730
rect 17618 8676 17642 8678
rect 17698 8676 17722 8678
rect 17778 8676 17802 8678
rect 17562 8656 17858 8676
rect 17972 8634 18000 8978
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 17972 8430 18000 8570
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 17132 7336 17184 7342
rect 17132 7278 17184 7284
rect 17144 6934 17172 7278
rect 17132 6928 17184 6934
rect 17132 6870 17184 6876
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 16500 5914 16528 6734
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 17144 5234 17172 6870
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 16488 5092 16540 5098
rect 16488 5034 16540 5040
rect 16500 4486 16528 5034
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16316 2746 16436 2774
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 16316 2310 16344 2746
rect 16500 2582 16528 4422
rect 17144 4146 17172 5170
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 17144 3670 17172 4082
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 17144 2922 17172 3606
rect 17236 2990 17264 8298
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 17328 7154 17356 7686
rect 17420 7342 17448 8026
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 17562 7644 17858 7664
rect 17618 7642 17642 7644
rect 17698 7642 17722 7644
rect 17778 7642 17802 7644
rect 17640 7590 17642 7642
rect 17704 7590 17716 7642
rect 17778 7590 17780 7642
rect 17618 7588 17642 7590
rect 17698 7588 17722 7590
rect 17778 7588 17802 7590
rect 17562 7568 17858 7588
rect 17408 7336 17460 7342
rect 17408 7278 17460 7284
rect 17328 7126 17448 7154
rect 17420 5778 17448 7126
rect 17972 7002 18000 7822
rect 18064 7206 18092 7890
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 17960 6996 18012 7002
rect 17960 6938 18012 6944
rect 18064 6866 18092 7142
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 17562 6556 17858 6576
rect 17618 6554 17642 6556
rect 17698 6554 17722 6556
rect 17778 6554 17802 6556
rect 17640 6502 17642 6554
rect 17704 6502 17716 6554
rect 17778 6502 17780 6554
rect 17618 6500 17642 6502
rect 17698 6500 17722 6502
rect 17778 6500 17802 6502
rect 17562 6480 17858 6500
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17420 5642 17540 5658
rect 17316 5636 17368 5642
rect 17316 5578 17368 5584
rect 17420 5636 17552 5642
rect 17420 5630 17500 5636
rect 17328 4826 17356 5578
rect 17420 5166 17448 5630
rect 17500 5578 17552 5584
rect 17562 5468 17858 5488
rect 17618 5466 17642 5468
rect 17698 5466 17722 5468
rect 17778 5466 17802 5468
rect 17640 5414 17642 5466
rect 17704 5414 17716 5466
rect 17778 5414 17780 5466
rect 17618 5412 17642 5414
rect 17698 5412 17722 5414
rect 17778 5412 17802 5414
rect 17562 5392 17858 5412
rect 17408 5160 17460 5166
rect 17408 5102 17460 5108
rect 17972 5030 18000 5714
rect 18156 5574 18184 10474
rect 18248 9178 18276 10542
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18340 8090 18368 10662
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 18524 10554 18552 11222
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 18432 10526 18552 10554
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 17316 4820 17368 4826
rect 17316 4762 17368 4768
rect 17972 4690 18000 4966
rect 17960 4684 18012 4690
rect 17960 4626 18012 4632
rect 17562 4380 17858 4400
rect 17618 4378 17642 4380
rect 17698 4378 17722 4380
rect 17778 4378 17802 4380
rect 17640 4326 17642 4378
rect 17704 4326 17716 4378
rect 17778 4326 17780 4378
rect 17618 4324 17642 4326
rect 17698 4324 17722 4326
rect 17778 4324 17802 4326
rect 17562 4304 17858 4324
rect 18156 3602 18184 5510
rect 18340 4690 18368 8026
rect 18432 6118 18460 10526
rect 18616 9518 18644 10610
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18708 6934 18736 8366
rect 18800 8362 18828 12038
rect 18984 11082 19012 13330
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19076 11694 19104 12038
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 19260 11150 19288 11834
rect 19996 11354 20024 12854
rect 20088 12434 20116 35022
rect 20996 34468 21048 34474
rect 20996 34410 21048 34416
rect 20720 34400 20772 34406
rect 20720 34342 20772 34348
rect 20732 34134 20760 34342
rect 20720 34128 20772 34134
rect 20720 34070 20772 34076
rect 21008 33998 21036 34410
rect 20996 33992 21048 33998
rect 20996 33934 21048 33940
rect 21640 33992 21692 33998
rect 21640 33934 21692 33940
rect 20720 33516 20772 33522
rect 20720 33458 20772 33464
rect 20260 32768 20312 32774
rect 20260 32710 20312 32716
rect 20444 32768 20496 32774
rect 20444 32710 20496 32716
rect 20168 32360 20220 32366
rect 20168 32302 20220 32308
rect 20180 32026 20208 32302
rect 20272 32026 20300 32710
rect 20456 32434 20484 32710
rect 20444 32428 20496 32434
rect 20444 32370 20496 32376
rect 20168 32020 20220 32026
rect 20168 31962 20220 31968
rect 20260 32020 20312 32026
rect 20260 31962 20312 31968
rect 20732 31754 20760 33458
rect 21008 32230 21036 33934
rect 21180 33856 21232 33862
rect 21180 33798 21232 33804
rect 21192 33522 21220 33798
rect 21652 33658 21680 33934
rect 21640 33652 21692 33658
rect 21640 33594 21692 33600
rect 21836 33590 21864 35090
rect 27080 34746 27108 35158
rect 29932 35154 29960 36853
rect 32692 35222 32720 36853
rect 32680 35216 32732 35222
rect 32680 35158 32732 35164
rect 34992 35154 35020 36853
rect 29920 35148 29972 35154
rect 29920 35090 29972 35096
rect 34980 35148 35032 35154
rect 34980 35090 35032 35096
rect 29276 35080 29328 35086
rect 29276 35022 29328 35028
rect 28632 34844 28928 34864
rect 28688 34842 28712 34844
rect 28768 34842 28792 34844
rect 28848 34842 28872 34844
rect 28710 34790 28712 34842
rect 28774 34790 28786 34842
rect 28848 34790 28850 34842
rect 28688 34788 28712 34790
rect 28768 34788 28792 34790
rect 28848 34788 28872 34790
rect 28632 34768 28928 34788
rect 27068 34740 27120 34746
rect 27068 34682 27120 34688
rect 23020 34536 23072 34542
rect 23020 34478 23072 34484
rect 21916 34400 21968 34406
rect 21916 34342 21968 34348
rect 21928 34134 21956 34342
rect 23032 34202 23060 34478
rect 23756 34400 23808 34406
rect 23756 34342 23808 34348
rect 23097 34300 23393 34320
rect 23153 34298 23177 34300
rect 23233 34298 23257 34300
rect 23313 34298 23337 34300
rect 23175 34246 23177 34298
rect 23239 34246 23251 34298
rect 23313 34246 23315 34298
rect 23153 34244 23177 34246
rect 23233 34244 23257 34246
rect 23313 34244 23337 34246
rect 23097 34224 23393 34244
rect 23768 34202 23796 34342
rect 23020 34196 23072 34202
rect 23020 34138 23072 34144
rect 23756 34196 23808 34202
rect 23756 34138 23808 34144
rect 21916 34128 21968 34134
rect 21916 34070 21968 34076
rect 21824 33584 21876 33590
rect 21824 33526 21876 33532
rect 21180 33516 21232 33522
rect 21180 33458 21232 33464
rect 21928 33386 21956 34070
rect 23572 34060 23624 34066
rect 23572 34002 23624 34008
rect 23584 33862 23612 34002
rect 23572 33856 23624 33862
rect 23572 33798 23624 33804
rect 21916 33380 21968 33386
rect 21916 33322 21968 33328
rect 21272 33312 21324 33318
rect 21272 33254 21324 33260
rect 21284 32910 21312 33254
rect 21272 32904 21324 32910
rect 21272 32846 21324 32852
rect 21284 32502 21312 32846
rect 21272 32496 21324 32502
rect 21272 32438 21324 32444
rect 21180 32292 21232 32298
rect 21180 32234 21232 32240
rect 20996 32224 21048 32230
rect 20996 32166 21048 32172
rect 20720 31748 20772 31754
rect 20720 31690 20772 31696
rect 20732 31482 20760 31690
rect 20720 31476 20772 31482
rect 20720 31418 20772 31424
rect 20536 30796 20588 30802
rect 20536 30738 20588 30744
rect 20352 30660 20404 30666
rect 20352 30602 20404 30608
rect 20364 30258 20392 30602
rect 20352 30252 20404 30258
rect 20352 30194 20404 30200
rect 20548 29510 20576 30738
rect 21088 30592 21140 30598
rect 21088 30534 21140 30540
rect 21100 30258 21128 30534
rect 21088 30252 21140 30258
rect 21088 30194 21140 30200
rect 20996 30184 21048 30190
rect 20916 30132 20996 30138
rect 20916 30126 21048 30132
rect 20916 30110 21036 30126
rect 20916 29646 20944 30110
rect 21192 30054 21220 32234
rect 21284 32026 21312 32438
rect 21928 32298 21956 33322
rect 23097 33212 23393 33232
rect 23153 33210 23177 33212
rect 23233 33210 23257 33212
rect 23313 33210 23337 33212
rect 23175 33158 23177 33210
rect 23239 33158 23251 33210
rect 23313 33158 23315 33210
rect 23153 33156 23177 33158
rect 23233 33156 23257 33158
rect 23313 33156 23337 33158
rect 23097 33136 23393 33156
rect 23584 33046 23612 33798
rect 23664 33312 23716 33318
rect 23664 33254 23716 33260
rect 23572 33040 23624 33046
rect 23572 32982 23624 32988
rect 22836 32904 22888 32910
rect 22836 32846 22888 32852
rect 21916 32292 21968 32298
rect 21916 32234 21968 32240
rect 21364 32224 21416 32230
rect 21364 32166 21416 32172
rect 21272 32020 21324 32026
rect 21272 31962 21324 31968
rect 21376 30190 21404 32166
rect 21928 31958 21956 32234
rect 22848 32230 22876 32846
rect 23676 32842 23704 33254
rect 23768 32978 23796 34138
rect 23940 33992 23992 33998
rect 23940 33934 23992 33940
rect 23756 32972 23808 32978
rect 23756 32914 23808 32920
rect 23664 32836 23716 32842
rect 23664 32778 23716 32784
rect 23480 32428 23532 32434
rect 23480 32370 23532 32376
rect 22100 32224 22152 32230
rect 22100 32166 22152 32172
rect 22836 32224 22888 32230
rect 22836 32166 22888 32172
rect 23020 32224 23072 32230
rect 23020 32166 23072 32172
rect 21916 31952 21968 31958
rect 21916 31894 21968 31900
rect 22112 31822 22140 32166
rect 23032 31890 23060 32166
rect 23097 32124 23393 32144
rect 23153 32122 23177 32124
rect 23233 32122 23257 32124
rect 23313 32122 23337 32124
rect 23175 32070 23177 32122
rect 23239 32070 23251 32122
rect 23313 32070 23315 32122
rect 23153 32068 23177 32070
rect 23233 32068 23257 32070
rect 23313 32068 23337 32070
rect 23097 32048 23393 32068
rect 23020 31884 23072 31890
rect 23020 31826 23072 31832
rect 22100 31816 22152 31822
rect 22100 31758 22152 31764
rect 21364 30184 21416 30190
rect 21364 30126 21416 30132
rect 21180 30048 21232 30054
rect 21180 29990 21232 29996
rect 21192 29850 21220 29990
rect 21180 29844 21232 29850
rect 21180 29786 21232 29792
rect 20904 29640 20956 29646
rect 20904 29582 20956 29588
rect 21456 29640 21508 29646
rect 21456 29582 21508 29588
rect 20536 29504 20588 29510
rect 20536 29446 20588 29452
rect 20548 29102 20576 29446
rect 20916 29306 20944 29582
rect 20904 29300 20956 29306
rect 20904 29242 20956 29248
rect 20444 29096 20496 29102
rect 20444 29038 20496 29044
rect 20536 29096 20588 29102
rect 20536 29038 20588 29044
rect 20352 28960 20404 28966
rect 20352 28902 20404 28908
rect 20260 28620 20312 28626
rect 20260 28562 20312 28568
rect 20272 28082 20300 28562
rect 20364 28558 20392 28902
rect 20352 28552 20404 28558
rect 20352 28494 20404 28500
rect 20456 28082 20484 29038
rect 20260 28076 20312 28082
rect 20260 28018 20312 28024
rect 20444 28076 20496 28082
rect 20444 28018 20496 28024
rect 20812 28008 20864 28014
rect 20812 27950 20864 27956
rect 20720 27940 20772 27946
rect 20720 27882 20772 27888
rect 20732 27606 20760 27882
rect 20720 27600 20772 27606
rect 20720 27542 20772 27548
rect 20168 27328 20220 27334
rect 20168 27270 20220 27276
rect 20180 27130 20208 27270
rect 20168 27124 20220 27130
rect 20168 27066 20220 27072
rect 20732 26994 20760 27542
rect 20824 27538 20852 27950
rect 20812 27532 20864 27538
rect 20812 27474 20864 27480
rect 20720 26988 20772 26994
rect 20720 26930 20772 26936
rect 20444 26784 20496 26790
rect 20444 26726 20496 26732
rect 20168 26580 20220 26586
rect 20168 26522 20220 26528
rect 20180 25770 20208 26522
rect 20456 25906 20484 26726
rect 20732 26042 20760 26930
rect 20916 26382 20944 29242
rect 21468 28762 21496 29582
rect 22008 29504 22060 29510
rect 22008 29446 22060 29452
rect 21456 28756 21508 28762
rect 21456 28698 21508 28704
rect 22020 28626 22048 29446
rect 20996 28620 21048 28626
rect 20996 28562 21048 28568
rect 22008 28620 22060 28626
rect 22008 28562 22060 28568
rect 21008 27674 21036 28562
rect 21088 28552 21140 28558
rect 21088 28494 21140 28500
rect 21100 28218 21128 28494
rect 21088 28212 21140 28218
rect 21088 28154 21140 28160
rect 21088 28008 21140 28014
rect 21088 27950 21140 27956
rect 20996 27668 21048 27674
rect 20996 27610 21048 27616
rect 21100 27538 21128 27950
rect 21180 27872 21232 27878
rect 21180 27814 21232 27820
rect 21088 27532 21140 27538
rect 21088 27474 21140 27480
rect 21192 26994 21220 27814
rect 22112 27674 22140 31758
rect 22836 31272 22888 31278
rect 22836 31214 22888 31220
rect 22848 30802 22876 31214
rect 23097 31036 23393 31056
rect 23153 31034 23177 31036
rect 23233 31034 23257 31036
rect 23313 31034 23337 31036
rect 23175 30982 23177 31034
rect 23239 30982 23251 31034
rect 23313 30982 23315 31034
rect 23153 30980 23177 30982
rect 23233 30980 23257 30982
rect 23313 30980 23337 30982
rect 23097 30960 23393 30980
rect 23492 30938 23520 32370
rect 23676 32366 23704 32778
rect 23664 32360 23716 32366
rect 23664 32302 23716 32308
rect 23768 32298 23796 32914
rect 23952 32434 23980 33934
rect 28632 33756 28928 33776
rect 28688 33754 28712 33756
rect 28768 33754 28792 33756
rect 28848 33754 28872 33756
rect 28710 33702 28712 33754
rect 28774 33702 28786 33754
rect 28848 33702 28850 33754
rect 28688 33700 28712 33702
rect 28768 33700 28792 33702
rect 28848 33700 28872 33702
rect 28632 33680 28928 33700
rect 29288 33454 29316 35022
rect 29460 34944 29512 34950
rect 29460 34886 29512 34892
rect 32312 34944 32364 34950
rect 32312 34886 32364 34892
rect 32496 34944 32548 34950
rect 32496 34886 32548 34892
rect 29472 34542 29500 34886
rect 29460 34536 29512 34542
rect 29460 34478 29512 34484
rect 25320 33448 25372 33454
rect 25320 33390 25372 33396
rect 27804 33448 27856 33454
rect 27804 33390 27856 33396
rect 29276 33448 29328 33454
rect 29276 33390 29328 33396
rect 24308 33380 24360 33386
rect 24308 33322 24360 33328
rect 23940 32428 23992 32434
rect 23940 32370 23992 32376
rect 23756 32292 23808 32298
rect 23756 32234 23808 32240
rect 23572 31816 23624 31822
rect 23572 31758 23624 31764
rect 23584 31346 23612 31758
rect 24320 31346 24348 33322
rect 25332 32502 25360 33390
rect 25320 32496 25372 32502
rect 25320 32438 25372 32444
rect 26608 32428 26660 32434
rect 26608 32370 26660 32376
rect 25872 32224 25924 32230
rect 25872 32166 25924 32172
rect 26240 32224 26292 32230
rect 26240 32166 26292 32172
rect 25884 31890 25912 32166
rect 25872 31884 25924 31890
rect 25872 31826 25924 31832
rect 23572 31340 23624 31346
rect 23572 31282 23624 31288
rect 24308 31340 24360 31346
rect 24308 31282 24360 31288
rect 23480 30932 23532 30938
rect 23480 30874 23532 30880
rect 22836 30796 22888 30802
rect 22836 30738 22888 30744
rect 23584 30394 23612 31282
rect 23940 31272 23992 31278
rect 23940 31214 23992 31220
rect 23952 30938 23980 31214
rect 23940 30932 23992 30938
rect 23940 30874 23992 30880
rect 23940 30796 23992 30802
rect 23940 30738 23992 30744
rect 23952 30394 23980 30738
rect 23572 30388 23624 30394
rect 23572 30330 23624 30336
rect 23940 30388 23992 30394
rect 23940 30330 23992 30336
rect 23480 30252 23532 30258
rect 23480 30194 23532 30200
rect 23097 29948 23393 29968
rect 23153 29946 23177 29948
rect 23233 29946 23257 29948
rect 23313 29946 23337 29948
rect 23175 29894 23177 29946
rect 23239 29894 23251 29946
rect 23313 29894 23315 29946
rect 23153 29892 23177 29894
rect 23233 29892 23257 29894
rect 23313 29892 23337 29894
rect 23097 29872 23393 29892
rect 22560 29028 22612 29034
rect 22560 28970 22612 28976
rect 22572 28626 22600 28970
rect 23097 28860 23393 28880
rect 23153 28858 23177 28860
rect 23233 28858 23257 28860
rect 23313 28858 23337 28860
rect 23175 28806 23177 28858
rect 23239 28806 23251 28858
rect 23313 28806 23315 28858
rect 23153 28804 23177 28806
rect 23233 28804 23257 28806
rect 23313 28804 23337 28806
rect 23097 28784 23393 28804
rect 23492 28762 23520 30194
rect 24320 30122 24348 31282
rect 25320 31136 25372 31142
rect 25320 31078 25372 31084
rect 25332 30938 25360 31078
rect 25320 30932 25372 30938
rect 25320 30874 25372 30880
rect 24860 30660 24912 30666
rect 24860 30602 24912 30608
rect 24768 30388 24820 30394
rect 24768 30330 24820 30336
rect 24308 30116 24360 30122
rect 24308 30058 24360 30064
rect 24780 29714 24808 30330
rect 24872 30190 24900 30602
rect 24860 30184 24912 30190
rect 24860 30126 24912 30132
rect 24768 29708 24820 29714
rect 24768 29650 24820 29656
rect 24860 29572 24912 29578
rect 24860 29514 24912 29520
rect 24584 29164 24636 29170
rect 24584 29106 24636 29112
rect 24308 28960 24360 28966
rect 24308 28902 24360 28908
rect 23480 28756 23532 28762
rect 23480 28698 23532 28704
rect 24320 28626 24348 28902
rect 22560 28620 22612 28626
rect 22560 28562 22612 28568
rect 24308 28620 24360 28626
rect 24308 28562 24360 28568
rect 22572 27946 22600 28562
rect 23940 28484 23992 28490
rect 23940 28426 23992 28432
rect 22836 28416 22888 28422
rect 22836 28358 22888 28364
rect 23952 28370 23980 28426
rect 24124 28416 24176 28422
rect 23952 28364 24124 28370
rect 23952 28358 24176 28364
rect 22560 27940 22612 27946
rect 22560 27882 22612 27888
rect 22100 27668 22152 27674
rect 22100 27610 22152 27616
rect 22112 27470 22140 27610
rect 22376 27532 22428 27538
rect 22376 27474 22428 27480
rect 22468 27532 22520 27538
rect 22468 27474 22520 27480
rect 22100 27464 22152 27470
rect 22100 27406 22152 27412
rect 22192 27124 22244 27130
rect 22192 27066 22244 27072
rect 21180 26988 21232 26994
rect 21180 26930 21232 26936
rect 22204 26926 22232 27066
rect 22192 26920 22244 26926
rect 22192 26862 22244 26868
rect 21088 26784 21140 26790
rect 21088 26726 21140 26732
rect 21100 26450 21128 26726
rect 21088 26444 21140 26450
rect 21088 26386 21140 26392
rect 20904 26376 20956 26382
rect 20904 26318 20956 26324
rect 20720 26036 20772 26042
rect 20720 25978 20772 25984
rect 20444 25900 20496 25906
rect 20444 25842 20496 25848
rect 20168 25764 20220 25770
rect 20168 25706 20220 25712
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20180 23526 20208 24754
rect 21088 24744 21140 24750
rect 21088 24686 21140 24692
rect 20444 24676 20496 24682
rect 20444 24618 20496 24624
rect 20456 24410 20484 24618
rect 20536 24608 20588 24614
rect 20536 24550 20588 24556
rect 20812 24608 20864 24614
rect 20812 24550 20864 24556
rect 20444 24404 20496 24410
rect 20444 24346 20496 24352
rect 20168 23520 20220 23526
rect 20168 23462 20220 23468
rect 20180 22030 20208 23462
rect 20456 23338 20484 24346
rect 20364 23310 20484 23338
rect 20364 22438 20392 23310
rect 20444 23180 20496 23186
rect 20444 23122 20496 23128
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 20168 22024 20220 22030
rect 20220 21984 20300 22012
rect 20168 21966 20220 21972
rect 20168 20800 20220 20806
rect 20168 20742 20220 20748
rect 20180 20602 20208 20742
rect 20168 20596 20220 20602
rect 20168 20538 20220 20544
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 20180 18834 20208 20198
rect 20272 19854 20300 21984
rect 20352 21004 20404 21010
rect 20352 20946 20404 20952
rect 20364 20058 20392 20946
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20260 19848 20312 19854
rect 20260 19790 20312 19796
rect 20168 18828 20220 18834
rect 20168 18770 20220 18776
rect 20272 18358 20300 19790
rect 20364 19310 20392 19994
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 20456 19174 20484 23122
rect 20548 22506 20576 24550
rect 20628 23588 20680 23594
rect 20628 23530 20680 23536
rect 20536 22500 20588 22506
rect 20536 22442 20588 22448
rect 20640 22438 20668 23530
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 20628 22432 20680 22438
rect 20628 22374 20680 22380
rect 20732 21690 20760 23122
rect 20824 23118 20852 24550
rect 21100 24410 21128 24686
rect 21088 24404 21140 24410
rect 21088 24346 21140 24352
rect 20996 24200 21048 24206
rect 20996 24142 21048 24148
rect 21364 24200 21416 24206
rect 21364 24142 21416 24148
rect 21008 23526 21036 24142
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 21376 23322 21404 24142
rect 21364 23316 21416 23322
rect 21364 23258 21416 23264
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 21732 23112 21784 23118
rect 21732 23054 21784 23060
rect 21456 22228 21508 22234
rect 21456 22170 21508 22176
rect 20720 21684 20772 21690
rect 20720 21626 20772 21632
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 21008 20398 21036 20878
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20626 19408 20682 19417
rect 20626 19343 20628 19352
rect 20680 19343 20682 19352
rect 20628 19314 20680 19320
rect 20732 19242 20760 19790
rect 20904 19372 20956 19378
rect 20824 19352 20904 19360
rect 20812 19346 20904 19352
rect 20864 19332 20904 19346
rect 20904 19314 20956 19320
rect 21008 19310 21036 20334
rect 21364 19984 21416 19990
rect 21284 19944 21364 19972
rect 20812 19288 20864 19294
rect 20996 19304 21048 19310
rect 20996 19246 21048 19252
rect 20720 19236 20772 19242
rect 20720 19178 20772 19184
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 20260 18352 20312 18358
rect 20260 18294 20312 18300
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20272 14550 20300 14758
rect 20260 14544 20312 14550
rect 20260 14486 20312 14492
rect 20088 12406 20208 12434
rect 20076 12368 20128 12374
rect 20076 12310 20128 12316
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 19800 11212 19852 11218
rect 19800 11154 19852 11160
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 18972 11076 19024 11082
rect 18972 11018 19024 11024
rect 19260 10606 19288 11086
rect 19812 10810 19840 11154
rect 19800 10804 19852 10810
rect 19800 10746 19852 10752
rect 19248 10600 19300 10606
rect 19248 10542 19300 10548
rect 19812 9518 19840 10746
rect 19996 10690 20024 11290
rect 19904 10662 20024 10690
rect 19800 9512 19852 9518
rect 19800 9454 19852 9460
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18892 7154 18920 8774
rect 18984 8430 19012 8774
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 19156 8356 19208 8362
rect 19156 8298 19208 8304
rect 18892 7126 19012 7154
rect 18696 6928 18748 6934
rect 18696 6870 18748 6876
rect 18984 6746 19012 7126
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 18708 6718 19012 6746
rect 18708 6662 18736 6718
rect 18984 6662 19012 6718
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18880 6656 18932 6662
rect 18880 6598 18932 6604
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 18892 6254 18920 6598
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18432 5778 18460 6054
rect 18420 5772 18472 5778
rect 18420 5714 18472 5720
rect 19076 5574 19104 6802
rect 19064 5568 19116 5574
rect 19064 5510 19116 5516
rect 19168 4690 19196 8298
rect 19616 7744 19668 7750
rect 19616 7686 19668 7692
rect 19628 7342 19656 7686
rect 19720 7546 19748 8910
rect 19800 8628 19852 8634
rect 19800 8570 19852 8576
rect 19708 7540 19760 7546
rect 19708 7482 19760 7488
rect 19812 7342 19840 8570
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19524 6928 19576 6934
rect 19524 6870 19576 6876
rect 19536 6322 19564 6870
rect 19628 6730 19656 7278
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 19628 5710 19656 6666
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 19904 4690 19932 10662
rect 19984 10532 20036 10538
rect 19984 10474 20036 10480
rect 19996 10266 20024 10474
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19984 10056 20036 10062
rect 19984 9998 20036 10004
rect 19996 9722 20024 9998
rect 19984 9716 20036 9722
rect 19984 9658 20036 9664
rect 20088 9450 20116 12310
rect 20180 12306 20208 12406
rect 20168 12300 20220 12306
rect 20168 12242 20220 12248
rect 20180 11898 20208 12242
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 20364 11218 20392 18702
rect 21284 18170 21312 19944
rect 21468 19972 21496 22170
rect 21744 22166 21772 23054
rect 21824 22704 21876 22710
rect 21824 22646 21876 22652
rect 21836 22166 21864 22646
rect 21732 22160 21784 22166
rect 21732 22102 21784 22108
rect 21824 22160 21876 22166
rect 21824 22102 21876 22108
rect 21824 21956 21876 21962
rect 21824 21898 21876 21904
rect 21836 21554 21864 21898
rect 21916 21888 21968 21894
rect 21916 21830 21968 21836
rect 21928 21690 21956 21830
rect 21916 21684 21968 21690
rect 21916 21626 21968 21632
rect 21928 21554 21956 21626
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 21916 21548 21968 21554
rect 21916 21490 21968 21496
rect 22204 20466 22232 26862
rect 22284 26444 22336 26450
rect 22284 26386 22336 26392
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 21416 19944 21496 19972
rect 21364 19926 21416 19932
rect 21640 19780 21692 19786
rect 21640 19722 21692 19728
rect 21652 19514 21680 19722
rect 22100 19712 22152 19718
rect 22100 19654 22152 19660
rect 21640 19508 21692 19514
rect 21640 19450 21692 19456
rect 22112 19310 22140 19654
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 21100 18154 21312 18170
rect 21088 18148 21312 18154
rect 21140 18142 21312 18148
rect 21364 18148 21416 18154
rect 21088 18090 21140 18096
rect 21364 18090 21416 18096
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 20444 16652 20496 16658
rect 20444 16594 20496 16600
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 20456 16454 20484 16594
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 20456 14958 20484 16390
rect 20640 16250 20668 16594
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20732 15978 20760 17682
rect 20904 17060 20956 17066
rect 20904 17002 20956 17008
rect 20812 16516 20864 16522
rect 20812 16458 20864 16464
rect 20536 15972 20588 15978
rect 20536 15914 20588 15920
rect 20720 15972 20772 15978
rect 20720 15914 20772 15920
rect 20548 15706 20576 15914
rect 20824 15910 20852 16458
rect 20916 16250 20944 17002
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20444 14952 20496 14958
rect 20444 14894 20496 14900
rect 20732 14890 20760 15642
rect 20720 14884 20772 14890
rect 20720 14826 20772 14832
rect 20732 14550 20760 14826
rect 20720 14544 20772 14550
rect 20720 14486 20772 14492
rect 20732 13530 20760 14486
rect 20824 13870 20852 15846
rect 20916 14618 20944 16186
rect 21008 16114 21036 16730
rect 21100 16590 21128 18090
rect 21272 18080 21324 18086
rect 21272 18022 21324 18028
rect 21284 17746 21312 18022
rect 21376 17882 21404 18090
rect 21364 17876 21416 17882
rect 21364 17818 21416 17824
rect 22100 17808 22152 17814
rect 22100 17750 22152 17756
rect 21272 17740 21324 17746
rect 21272 17682 21324 17688
rect 22112 17134 22140 17750
rect 22100 17128 22152 17134
rect 22100 17070 22152 17076
rect 22112 16658 22140 17070
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 21916 16584 21968 16590
rect 21916 16526 21968 16532
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 21732 16108 21784 16114
rect 21732 16050 21784 16056
rect 21744 15570 21772 16050
rect 21928 15706 21956 16526
rect 22008 15904 22060 15910
rect 22008 15846 22060 15852
rect 21916 15700 21968 15706
rect 21916 15642 21968 15648
rect 22020 15638 22048 15846
rect 22008 15632 22060 15638
rect 22008 15574 22060 15580
rect 21732 15564 21784 15570
rect 21732 15506 21784 15512
rect 22296 15178 22324 26386
rect 22388 26382 22416 27474
rect 22376 26376 22428 26382
rect 22376 26318 22428 26324
rect 22480 26042 22508 27474
rect 22468 26036 22520 26042
rect 22468 25978 22520 25984
rect 22572 24614 22600 27882
rect 22848 27878 22876 28358
rect 23952 28342 24164 28358
rect 23952 28098 23980 28342
rect 23952 28070 24072 28098
rect 24044 28014 24072 28070
rect 24032 28008 24084 28014
rect 24032 27950 24084 27956
rect 22836 27872 22888 27878
rect 22836 27814 22888 27820
rect 23572 27872 23624 27878
rect 23572 27814 23624 27820
rect 22652 27328 22704 27334
rect 22652 27270 22704 27276
rect 22744 27328 22796 27334
rect 22744 27270 22796 27276
rect 22664 26926 22692 27270
rect 22756 26994 22784 27270
rect 22848 27130 22876 27814
rect 23097 27772 23393 27792
rect 23153 27770 23177 27772
rect 23233 27770 23257 27772
rect 23313 27770 23337 27772
rect 23175 27718 23177 27770
rect 23239 27718 23251 27770
rect 23313 27718 23315 27770
rect 23153 27716 23177 27718
rect 23233 27716 23257 27718
rect 23313 27716 23337 27718
rect 23097 27696 23393 27716
rect 22836 27124 22888 27130
rect 22836 27066 22888 27072
rect 22928 27056 22980 27062
rect 22928 26998 22980 27004
rect 22744 26988 22796 26994
rect 22744 26930 22796 26936
rect 22652 26920 22704 26926
rect 22652 26862 22704 26868
rect 22940 26586 22968 26998
rect 23020 26920 23072 26926
rect 23020 26862 23072 26868
rect 22928 26580 22980 26586
rect 22928 26522 22980 26528
rect 22940 25362 22968 26522
rect 23032 26518 23060 26862
rect 23097 26684 23393 26704
rect 23153 26682 23177 26684
rect 23233 26682 23257 26684
rect 23313 26682 23337 26684
rect 23175 26630 23177 26682
rect 23239 26630 23251 26682
rect 23313 26630 23315 26682
rect 23153 26628 23177 26630
rect 23233 26628 23257 26630
rect 23313 26628 23337 26630
rect 23097 26608 23393 26628
rect 23020 26512 23072 26518
rect 23020 26454 23072 26460
rect 23032 25838 23060 26454
rect 23020 25832 23072 25838
rect 23020 25774 23072 25780
rect 23480 25832 23532 25838
rect 23480 25774 23532 25780
rect 23097 25596 23393 25616
rect 23153 25594 23177 25596
rect 23233 25594 23257 25596
rect 23313 25594 23337 25596
rect 23175 25542 23177 25594
rect 23239 25542 23251 25594
rect 23313 25542 23315 25594
rect 23153 25540 23177 25542
rect 23233 25540 23257 25542
rect 23313 25540 23337 25542
rect 23097 25520 23393 25540
rect 23492 25362 23520 25774
rect 22928 25356 22980 25362
rect 22928 25298 22980 25304
rect 23480 25356 23532 25362
rect 23480 25298 23532 25304
rect 22940 24818 22968 25298
rect 22928 24812 22980 24818
rect 22928 24754 22980 24760
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 22560 24608 22612 24614
rect 22560 24550 22612 24556
rect 22376 24336 22428 24342
rect 22376 24278 22428 24284
rect 22388 23186 22416 24278
rect 22376 23180 22428 23186
rect 22376 23122 22428 23128
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22388 21690 22416 21966
rect 22376 21684 22428 21690
rect 22376 21626 22428 21632
rect 22572 21536 22600 24550
rect 22940 24410 22968 24754
rect 23020 24676 23072 24682
rect 23020 24618 23072 24624
rect 22928 24404 22980 24410
rect 22928 24346 22980 24352
rect 23032 24342 23060 24618
rect 23097 24508 23393 24528
rect 23153 24506 23177 24508
rect 23233 24506 23257 24508
rect 23313 24506 23337 24508
rect 23175 24454 23177 24506
rect 23239 24454 23251 24506
rect 23313 24454 23315 24506
rect 23153 24452 23177 24454
rect 23233 24452 23257 24454
rect 23313 24452 23337 24454
rect 23097 24432 23393 24452
rect 23020 24336 23072 24342
rect 23020 24278 23072 24284
rect 23020 24064 23072 24070
rect 23020 24006 23072 24012
rect 23032 23254 23060 24006
rect 23492 23662 23520 24754
rect 23480 23656 23532 23662
rect 23480 23598 23532 23604
rect 23097 23420 23393 23440
rect 23153 23418 23177 23420
rect 23233 23418 23257 23420
rect 23313 23418 23337 23420
rect 23175 23366 23177 23418
rect 23239 23366 23251 23418
rect 23313 23366 23315 23418
rect 23153 23364 23177 23366
rect 23233 23364 23257 23366
rect 23313 23364 23337 23366
rect 23097 23344 23393 23364
rect 23492 23254 23520 23598
rect 23584 23594 23612 27814
rect 24596 27402 24624 29106
rect 24768 28688 24820 28694
rect 24768 28630 24820 28636
rect 24780 28014 24808 28630
rect 24872 28082 24900 29514
rect 25136 29504 25188 29510
rect 25136 29446 25188 29452
rect 25148 29034 25176 29446
rect 25332 29306 25360 30874
rect 26252 30734 26280 32166
rect 26516 32020 26568 32026
rect 26516 31962 26568 31968
rect 26528 31210 26556 31962
rect 26516 31204 26568 31210
rect 26516 31146 26568 31152
rect 26528 30870 26556 31146
rect 26516 30864 26568 30870
rect 26516 30806 26568 30812
rect 26240 30728 26292 30734
rect 26240 30670 26292 30676
rect 26252 30190 26280 30670
rect 26148 30184 26200 30190
rect 26148 30126 26200 30132
rect 26240 30184 26292 30190
rect 26240 30126 26292 30132
rect 25872 30048 25924 30054
rect 25872 29990 25924 29996
rect 25504 29708 25556 29714
rect 25504 29650 25556 29656
rect 25516 29306 25544 29650
rect 25320 29300 25372 29306
rect 25320 29242 25372 29248
rect 25504 29300 25556 29306
rect 25504 29242 25556 29248
rect 25136 29028 25188 29034
rect 25136 28970 25188 28976
rect 25332 28762 25360 29242
rect 25596 28960 25648 28966
rect 25596 28902 25648 28908
rect 25320 28756 25372 28762
rect 25320 28698 25372 28704
rect 25228 28416 25280 28422
rect 25228 28358 25280 28364
rect 24860 28076 24912 28082
rect 24860 28018 24912 28024
rect 24768 28008 24820 28014
rect 24768 27950 24820 27956
rect 24032 27396 24084 27402
rect 24032 27338 24084 27344
rect 24584 27396 24636 27402
rect 24584 27338 24636 27344
rect 24044 26926 24072 27338
rect 24780 27130 24808 27950
rect 25240 27674 25268 28358
rect 25332 28014 25360 28698
rect 25320 28008 25372 28014
rect 25320 27950 25372 27956
rect 25228 27668 25280 27674
rect 25228 27610 25280 27616
rect 25044 27532 25096 27538
rect 25044 27474 25096 27480
rect 25136 27532 25188 27538
rect 25136 27474 25188 27480
rect 24768 27124 24820 27130
rect 24768 27066 24820 27072
rect 25056 27062 25084 27474
rect 25044 27056 25096 27062
rect 25044 26998 25096 27004
rect 24032 26920 24084 26926
rect 24032 26862 24084 26868
rect 24860 26852 24912 26858
rect 24860 26794 24912 26800
rect 24872 26382 24900 26794
rect 24952 26784 25004 26790
rect 24952 26726 25004 26732
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 24964 26314 24992 26726
rect 24952 26308 25004 26314
rect 24952 26250 25004 26256
rect 24964 25770 24992 26250
rect 23848 25764 23900 25770
rect 23848 25706 23900 25712
rect 24124 25764 24176 25770
rect 24124 25706 24176 25712
rect 24952 25764 25004 25770
rect 24952 25706 25004 25712
rect 23860 25158 23888 25706
rect 23940 25696 23992 25702
rect 23940 25638 23992 25644
rect 23952 25430 23980 25638
rect 23940 25424 23992 25430
rect 23940 25366 23992 25372
rect 23848 25152 23900 25158
rect 23848 25094 23900 25100
rect 23756 24744 23808 24750
rect 23756 24686 23808 24692
rect 23664 24064 23716 24070
rect 23664 24006 23716 24012
rect 23572 23588 23624 23594
rect 23572 23530 23624 23536
rect 23020 23248 23072 23254
rect 23020 23190 23072 23196
rect 23480 23248 23532 23254
rect 23480 23190 23532 23196
rect 23032 22574 23060 23190
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23020 22568 23072 22574
rect 23020 22510 23072 22516
rect 23097 22332 23393 22352
rect 23153 22330 23177 22332
rect 23233 22330 23257 22332
rect 23313 22330 23337 22332
rect 23175 22278 23177 22330
rect 23239 22278 23251 22330
rect 23313 22278 23315 22330
rect 23153 22276 23177 22278
rect 23233 22276 23257 22278
rect 23313 22276 23337 22278
rect 23097 22256 23393 22276
rect 22744 22092 22796 22098
rect 22744 22034 22796 22040
rect 22652 21548 22704 21554
rect 22388 21508 22652 21536
rect 22388 21010 22416 21508
rect 22652 21490 22704 21496
rect 22468 21412 22520 21418
rect 22468 21354 22520 21360
rect 22480 21078 22508 21354
rect 22468 21072 22520 21078
rect 22468 21014 22520 21020
rect 22756 21010 22784 22034
rect 22928 21480 22980 21486
rect 22928 21422 22980 21428
rect 22940 21350 22968 21422
rect 23032 21418 23152 21434
rect 23032 21412 23164 21418
rect 23032 21406 23112 21412
rect 22928 21344 22980 21350
rect 22928 21286 22980 21292
rect 22376 21004 22428 21010
rect 22376 20946 22428 20952
rect 22744 21004 22796 21010
rect 22744 20946 22796 20952
rect 22560 20460 22612 20466
rect 22560 20402 22612 20408
rect 22480 19417 22508 19443
rect 22466 19408 22522 19417
rect 22466 19343 22468 19352
rect 22520 19343 22522 19352
rect 22468 19314 22520 19320
rect 22480 16250 22508 19314
rect 22572 19242 22600 20402
rect 23032 20398 23060 21406
rect 23112 21354 23164 21360
rect 23097 21244 23393 21264
rect 23153 21242 23177 21244
rect 23233 21242 23257 21244
rect 23313 21242 23337 21244
rect 23175 21190 23177 21242
rect 23239 21190 23251 21242
rect 23313 21190 23315 21242
rect 23153 21188 23177 21190
rect 23233 21188 23257 21190
rect 23313 21188 23337 21190
rect 23097 21168 23393 21188
rect 23492 20398 23520 22918
rect 23572 22704 23624 22710
rect 23572 22646 23624 22652
rect 23584 22098 23612 22646
rect 23676 22574 23704 24006
rect 23664 22568 23716 22574
rect 23664 22510 23716 22516
rect 23572 22092 23624 22098
rect 23572 22034 23624 22040
rect 23584 21486 23612 22034
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 23768 21162 23796 24686
rect 23860 24682 23888 25094
rect 23952 24750 23980 25366
rect 24136 25362 24164 25706
rect 24124 25356 24176 25362
rect 24124 25298 24176 25304
rect 25056 24750 25084 26998
rect 23940 24744 23992 24750
rect 23940 24686 23992 24692
rect 25044 24744 25096 24750
rect 25044 24686 25096 24692
rect 23848 24676 23900 24682
rect 23848 24618 23900 24624
rect 23860 24274 23888 24618
rect 23952 24342 23980 24686
rect 25148 24410 25176 27474
rect 25320 26988 25372 26994
rect 25320 26930 25372 26936
rect 25332 26586 25360 26930
rect 25320 26580 25372 26586
rect 25320 26522 25372 26528
rect 25332 26450 25360 26522
rect 25320 26444 25372 26450
rect 25320 26386 25372 26392
rect 25412 26444 25464 26450
rect 25412 26386 25464 26392
rect 25320 25832 25372 25838
rect 25424 25820 25452 26386
rect 25504 26308 25556 26314
rect 25504 26250 25556 26256
rect 25372 25792 25452 25820
rect 25320 25774 25372 25780
rect 25332 25498 25360 25774
rect 25320 25492 25372 25498
rect 25320 25434 25372 25440
rect 25228 24608 25280 24614
rect 25228 24550 25280 24556
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 23940 24336 23992 24342
rect 23940 24278 23992 24284
rect 23848 24268 23900 24274
rect 23848 24210 23900 24216
rect 24400 24064 24452 24070
rect 24400 24006 24452 24012
rect 24412 23662 24440 24006
rect 23848 23656 23900 23662
rect 23848 23598 23900 23604
rect 24400 23656 24452 23662
rect 24400 23598 24452 23604
rect 23860 23050 23888 23598
rect 24308 23588 24360 23594
rect 24308 23530 24360 23536
rect 23848 23044 23900 23050
rect 23848 22986 23900 22992
rect 23848 22568 23900 22574
rect 23848 22510 23900 22516
rect 24032 22568 24084 22574
rect 24032 22510 24084 22516
rect 23860 21690 23888 22510
rect 23940 22432 23992 22438
rect 23940 22374 23992 22380
rect 23952 22030 23980 22374
rect 23940 22024 23992 22030
rect 23940 21966 23992 21972
rect 23848 21684 23900 21690
rect 23848 21626 23900 21632
rect 23940 21344 23992 21350
rect 23940 21286 23992 21292
rect 23768 21134 23888 21162
rect 23756 21004 23808 21010
rect 23756 20946 23808 20952
rect 23768 20398 23796 20946
rect 23860 20602 23888 21134
rect 23952 21010 23980 21286
rect 24044 21078 24072 22510
rect 24320 22094 24348 23530
rect 24412 23254 24440 23598
rect 24492 23588 24544 23594
rect 24492 23530 24544 23536
rect 24400 23248 24452 23254
rect 24400 23190 24452 23196
rect 24504 23100 24532 23530
rect 25148 23254 25176 24346
rect 25240 23730 25268 24550
rect 25516 24274 25544 26250
rect 25504 24268 25556 24274
rect 25504 24210 25556 24216
rect 25228 23724 25280 23730
rect 25228 23666 25280 23672
rect 25504 23588 25556 23594
rect 25504 23530 25556 23536
rect 25516 23322 25544 23530
rect 25504 23316 25556 23322
rect 25504 23258 25556 23264
rect 25136 23248 25188 23254
rect 25136 23190 25188 23196
rect 24768 23180 24820 23186
rect 24768 23122 24820 23128
rect 24412 23072 24532 23100
rect 24412 22574 24440 23072
rect 24780 22642 24808 23122
rect 24768 22636 24820 22642
rect 24768 22578 24820 22584
rect 24400 22568 24452 22574
rect 24400 22510 24452 22516
rect 24400 22094 24452 22098
rect 24320 22092 24452 22094
rect 24320 22066 24400 22092
rect 25608 22094 25636 28902
rect 25780 28552 25832 28558
rect 25780 28494 25832 28500
rect 25688 28416 25740 28422
rect 25688 28358 25740 28364
rect 25700 28150 25728 28358
rect 25792 28218 25820 28494
rect 25780 28212 25832 28218
rect 25780 28154 25832 28160
rect 25688 28144 25740 28150
rect 25884 28098 25912 29990
rect 26160 29594 26188 30126
rect 26252 29714 26280 30126
rect 26424 30048 26476 30054
rect 26424 29990 26476 29996
rect 26436 29782 26464 29990
rect 26424 29776 26476 29782
rect 26424 29718 26476 29724
rect 26240 29708 26292 29714
rect 26240 29650 26292 29656
rect 26160 29578 26280 29594
rect 26160 29572 26292 29578
rect 26160 29566 26240 29572
rect 26240 29514 26292 29520
rect 25688 28086 25740 28092
rect 25792 28070 25912 28098
rect 25792 27878 25820 28070
rect 26056 27940 26108 27946
rect 26056 27882 26108 27888
rect 25780 27872 25832 27878
rect 25780 27814 25832 27820
rect 25792 23118 25820 27814
rect 25964 25764 26016 25770
rect 25964 25706 26016 25712
rect 25872 25696 25924 25702
rect 25872 25638 25924 25644
rect 25884 25430 25912 25638
rect 25872 25424 25924 25430
rect 25872 25366 25924 25372
rect 25976 24274 26004 25706
rect 25872 24268 25924 24274
rect 25872 24210 25924 24216
rect 25964 24268 26016 24274
rect 25964 24210 26016 24216
rect 25884 23202 25912 24210
rect 25884 23186 26004 23202
rect 25884 23180 26016 23186
rect 25884 23174 25964 23180
rect 25964 23122 26016 23128
rect 25780 23112 25832 23118
rect 25780 23054 25832 23060
rect 25780 22094 25832 22098
rect 25608 22092 25832 22094
rect 25608 22066 25780 22092
rect 24400 22034 24452 22040
rect 25700 22052 25780 22066
rect 24492 22024 24544 22030
rect 24492 21966 24544 21972
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 24504 21690 24532 21966
rect 24492 21684 24544 21690
rect 24492 21626 24544 21632
rect 24780 21622 24808 21966
rect 25504 21684 25556 21690
rect 25504 21626 25556 21632
rect 24768 21616 24820 21622
rect 24768 21558 24820 21564
rect 24860 21480 24912 21486
rect 24860 21422 24912 21428
rect 24872 21078 24900 21422
rect 25320 21412 25372 21418
rect 25320 21354 25372 21360
rect 24032 21072 24084 21078
rect 24032 21014 24084 21020
rect 24860 21072 24912 21078
rect 24860 21014 24912 21020
rect 23940 21004 23992 21010
rect 23940 20946 23992 20952
rect 23940 20800 23992 20806
rect 23940 20742 23992 20748
rect 23848 20596 23900 20602
rect 23848 20538 23900 20544
rect 23952 20466 23980 20742
rect 23940 20460 23992 20466
rect 23940 20402 23992 20408
rect 23020 20392 23072 20398
rect 23020 20334 23072 20340
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23756 20392 23808 20398
rect 23756 20334 23808 20340
rect 22836 20324 22888 20330
rect 22836 20266 22888 20272
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 22664 19310 22692 19654
rect 22652 19304 22704 19310
rect 22652 19246 22704 19252
rect 22744 19304 22796 19310
rect 22744 19246 22796 19252
rect 22560 19236 22612 19242
rect 22560 19178 22612 19184
rect 22652 18420 22704 18426
rect 22652 18362 22704 18368
rect 22664 17746 22692 18362
rect 22756 18290 22784 19246
rect 22744 18284 22796 18290
rect 22744 18226 22796 18232
rect 22848 17746 22876 20266
rect 23032 19922 23060 20334
rect 24044 20330 24072 21014
rect 25332 20942 25360 21354
rect 25516 21010 25544 21626
rect 25504 21004 25556 21010
rect 25504 20946 25556 20952
rect 25228 20936 25280 20942
rect 25228 20878 25280 20884
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 24768 20596 24820 20602
rect 24768 20538 24820 20544
rect 24032 20324 24084 20330
rect 24032 20266 24084 20272
rect 23572 20256 23624 20262
rect 23572 20198 23624 20204
rect 23097 20156 23393 20176
rect 23153 20154 23177 20156
rect 23233 20154 23257 20156
rect 23313 20154 23337 20156
rect 23175 20102 23177 20154
rect 23239 20102 23251 20154
rect 23313 20102 23315 20154
rect 23153 20100 23177 20102
rect 23233 20100 23257 20102
rect 23313 20100 23337 20102
rect 23097 20080 23393 20100
rect 23020 19916 23072 19922
rect 23020 19858 23072 19864
rect 23584 19378 23612 20198
rect 24780 19922 24808 20538
rect 24308 19916 24360 19922
rect 24308 19858 24360 19864
rect 24768 19916 24820 19922
rect 24768 19858 24820 19864
rect 24320 19514 24348 19858
rect 24308 19508 24360 19514
rect 24308 19450 24360 19456
rect 23572 19372 23624 19378
rect 23572 19314 23624 19320
rect 23020 19236 23072 19242
rect 23020 19178 23072 19184
rect 23664 19236 23716 19242
rect 23664 19178 23716 19184
rect 22652 17740 22704 17746
rect 22652 17682 22704 17688
rect 22836 17740 22888 17746
rect 22836 17682 22888 17688
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 22468 16244 22520 16250
rect 22468 16186 22520 16192
rect 21824 15156 21876 15162
rect 22296 15150 22416 15178
rect 21824 15098 21876 15104
rect 21732 14952 21784 14958
rect 21732 14894 21784 14900
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 20904 14612 20956 14618
rect 20904 14554 20956 14560
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20916 13802 20944 14554
rect 20904 13796 20956 13802
rect 20904 13738 20956 13744
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20732 12918 20760 13466
rect 20916 13190 20944 13738
rect 20996 13728 21048 13734
rect 20996 13670 21048 13676
rect 21008 13326 21036 13670
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 20904 13184 20956 13190
rect 20904 13126 20956 13132
rect 20916 12986 20944 13126
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 20720 12912 20772 12918
rect 20720 12854 20772 12860
rect 20444 12164 20496 12170
rect 20444 12106 20496 12112
rect 20456 11898 20484 12106
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 21284 11626 21312 12922
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21272 11620 21324 11626
rect 21272 11562 21324 11568
rect 20352 11212 20404 11218
rect 20352 11154 20404 11160
rect 20364 9518 20392 11154
rect 21284 10674 21312 11562
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 21376 10554 21404 12038
rect 21284 10526 21404 10554
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20824 10130 20852 10406
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20536 10056 20588 10062
rect 20536 9998 20588 10004
rect 20352 9512 20404 9518
rect 20352 9454 20404 9460
rect 20076 9444 20128 9450
rect 20076 9386 20128 9392
rect 20364 9178 20392 9454
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20168 8900 20220 8906
rect 20168 8842 20220 8848
rect 20180 8634 20208 8842
rect 20168 8628 20220 8634
rect 20168 8570 20220 8576
rect 20364 7954 20392 9114
rect 20548 8906 20576 9998
rect 21180 9648 21232 9654
rect 21180 9590 21232 9596
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 20536 8900 20588 8906
rect 20536 8842 20588 8848
rect 20352 7948 20404 7954
rect 20352 7890 20404 7896
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 20352 6792 20404 6798
rect 20352 6734 20404 6740
rect 20088 5914 20116 6734
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20272 6254 20300 6598
rect 20260 6248 20312 6254
rect 20260 6190 20312 6196
rect 20364 5914 20392 6734
rect 20076 5908 20128 5914
rect 20076 5850 20128 5856
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 20548 5370 20576 8842
rect 20640 8498 20668 9318
rect 20824 9042 20852 9318
rect 20916 9110 20944 9318
rect 20904 9104 20956 9110
rect 20904 9046 20956 9052
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 21192 8906 21220 9590
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 19156 4684 19208 4690
rect 19156 4626 19208 4632
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 20168 4684 20220 4690
rect 20168 4626 20220 4632
rect 18972 4480 19024 4486
rect 18972 4422 19024 4428
rect 18984 4078 19012 4422
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 19168 3602 19196 4626
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 19156 3596 19208 3602
rect 19156 3538 19208 3544
rect 17420 3194 17448 3538
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 17562 3292 17858 3312
rect 17618 3290 17642 3292
rect 17698 3290 17722 3292
rect 17778 3290 17802 3292
rect 17640 3238 17642 3290
rect 17704 3238 17716 3290
rect 17778 3238 17780 3290
rect 17618 3236 17642 3238
rect 17698 3236 17722 3238
rect 17778 3236 17802 3238
rect 17562 3216 17858 3236
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 17132 2916 17184 2922
rect 17132 2858 17184 2864
rect 17604 2650 17632 2994
rect 18340 2990 18368 3334
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18432 2650 18460 3470
rect 19168 3194 19196 3538
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 19904 2922 19932 4626
rect 20180 3942 20208 4626
rect 20640 4554 20668 8434
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 21100 6458 21128 7822
rect 21192 7546 21220 8842
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21284 6866 21312 10526
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 21376 9722 21404 10066
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21364 7336 21416 7342
rect 21468 7324 21496 14758
rect 21744 14618 21772 14894
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 21836 14074 21864 15098
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22296 14618 22324 14962
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 22296 13938 22324 14418
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 21732 13864 21784 13870
rect 21732 13806 21784 13812
rect 21744 13190 21772 13806
rect 21732 13184 21784 13190
rect 21732 13126 21784 13132
rect 21744 11218 21772 13126
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 21928 12442 21956 12922
rect 22008 12912 22060 12918
rect 22008 12854 22060 12860
rect 21916 12436 21968 12442
rect 21916 12378 21968 12384
rect 22020 12374 22048 12854
rect 22388 12714 22416 15150
rect 22480 15094 22508 16186
rect 22756 15978 22784 17478
rect 23032 16046 23060 19178
rect 23097 19068 23393 19088
rect 23153 19066 23177 19068
rect 23233 19066 23257 19068
rect 23313 19066 23337 19068
rect 23175 19014 23177 19066
rect 23239 19014 23251 19066
rect 23313 19014 23315 19066
rect 23153 19012 23177 19014
rect 23233 19012 23257 19014
rect 23313 19012 23337 19014
rect 23097 18992 23393 19012
rect 23676 18154 23704 19178
rect 23664 18148 23716 18154
rect 23664 18090 23716 18096
rect 24124 18148 24176 18154
rect 24124 18090 24176 18096
rect 23097 17980 23393 18000
rect 23153 17978 23177 17980
rect 23233 17978 23257 17980
rect 23313 17978 23337 17980
rect 23175 17926 23177 17978
rect 23239 17926 23251 17978
rect 23313 17926 23315 17978
rect 23153 17924 23177 17926
rect 23233 17924 23257 17926
rect 23313 17924 23337 17926
rect 23097 17904 23393 17924
rect 23676 17066 23704 18090
rect 24136 17882 24164 18090
rect 24124 17876 24176 17882
rect 24124 17818 24176 17824
rect 24584 17196 24636 17202
rect 24584 17138 24636 17144
rect 23664 17060 23716 17066
rect 23664 17002 23716 17008
rect 23097 16892 23393 16912
rect 23153 16890 23177 16892
rect 23233 16890 23257 16892
rect 23313 16890 23337 16892
rect 23175 16838 23177 16890
rect 23239 16838 23251 16890
rect 23313 16838 23315 16890
rect 23153 16836 23177 16838
rect 23233 16836 23257 16838
rect 23313 16836 23337 16838
rect 23097 16816 23393 16836
rect 23676 16658 23704 17002
rect 24596 16998 24624 17138
rect 23756 16992 23808 16998
rect 23756 16934 23808 16940
rect 24584 16992 24636 16998
rect 24584 16934 24636 16940
rect 23664 16652 23716 16658
rect 23664 16594 23716 16600
rect 23768 16538 23796 16934
rect 23676 16510 23796 16538
rect 24780 16522 24808 19858
rect 25136 19236 25188 19242
rect 25136 19178 25188 19184
rect 25148 18970 25176 19178
rect 25240 19174 25268 20878
rect 25332 20398 25360 20878
rect 25320 20392 25372 20398
rect 25320 20334 25372 20340
rect 25332 19990 25360 20334
rect 25596 20256 25648 20262
rect 25596 20198 25648 20204
rect 25320 19984 25372 19990
rect 25320 19926 25372 19932
rect 25332 19310 25360 19926
rect 25320 19304 25372 19310
rect 25320 19246 25372 19252
rect 25228 19168 25280 19174
rect 25228 19110 25280 19116
rect 25136 18964 25188 18970
rect 25136 18906 25188 18912
rect 25608 18873 25636 20198
rect 25700 19854 25728 22052
rect 25780 22034 25832 22040
rect 25976 20602 26004 23122
rect 26068 20602 26096 27882
rect 26252 27826 26280 29514
rect 26436 28914 26464 29718
rect 26344 28886 26464 28914
rect 26344 28762 26372 28886
rect 26332 28756 26384 28762
rect 26332 28698 26384 28704
rect 26344 28014 26372 28698
rect 26528 28694 26556 30806
rect 26620 30258 26648 32370
rect 27816 32366 27844 33390
rect 28172 33380 28224 33386
rect 28172 33322 28224 33328
rect 28184 32502 28212 33322
rect 28632 32668 28928 32688
rect 28688 32666 28712 32668
rect 28768 32666 28792 32668
rect 28848 32666 28872 32668
rect 28710 32614 28712 32666
rect 28774 32614 28786 32666
rect 28848 32614 28850 32666
rect 28688 32612 28712 32614
rect 28768 32612 28792 32614
rect 28848 32612 28872 32614
rect 28632 32592 28928 32612
rect 28172 32496 28224 32502
rect 28172 32438 28224 32444
rect 27804 32360 27856 32366
rect 29288 32314 29316 33390
rect 30012 33380 30064 33386
rect 30012 33322 30064 33328
rect 29460 32428 29512 32434
rect 29460 32370 29512 32376
rect 27804 32302 27856 32308
rect 26700 32292 26752 32298
rect 26700 32234 26752 32240
rect 26712 32026 26740 32234
rect 26700 32020 26752 32026
rect 26700 31962 26752 31968
rect 26608 30252 26660 30258
rect 26608 30194 26660 30200
rect 26516 28688 26568 28694
rect 26516 28630 26568 28636
rect 26332 28008 26384 28014
rect 26332 27950 26384 27956
rect 26608 28008 26660 28014
rect 26608 27950 26660 27956
rect 26252 27798 26464 27826
rect 26240 27532 26292 27538
rect 26240 27474 26292 27480
rect 26252 26926 26280 27474
rect 26332 27396 26384 27402
rect 26332 27338 26384 27344
rect 26240 26920 26292 26926
rect 26240 26862 26292 26868
rect 26344 26518 26372 27338
rect 26332 26512 26384 26518
rect 26332 26454 26384 26460
rect 26344 25906 26372 26454
rect 26332 25900 26384 25906
rect 26332 25842 26384 25848
rect 26436 24682 26464 27798
rect 26516 26036 26568 26042
rect 26516 25978 26568 25984
rect 26528 25906 26556 25978
rect 26516 25900 26568 25906
rect 26516 25842 26568 25848
rect 26424 24676 26476 24682
rect 26424 24618 26476 24624
rect 26148 22432 26200 22438
rect 26148 22374 26200 22380
rect 26160 22098 26188 22374
rect 26148 22092 26200 22098
rect 26148 22034 26200 22040
rect 26160 21350 26188 22034
rect 26436 21418 26464 24618
rect 26516 21888 26568 21894
rect 26516 21830 26568 21836
rect 26424 21412 26476 21418
rect 26424 21354 26476 21360
rect 26148 21344 26200 21350
rect 26148 21286 26200 21292
rect 26148 21004 26200 21010
rect 26148 20946 26200 20952
rect 25964 20596 26016 20602
rect 25964 20538 26016 20544
rect 26056 20596 26108 20602
rect 26056 20538 26108 20544
rect 25780 20392 25832 20398
rect 25780 20334 25832 20340
rect 25792 19922 25820 20334
rect 25780 19916 25832 19922
rect 25780 19858 25832 19864
rect 25688 19848 25740 19854
rect 25688 19790 25740 19796
rect 25688 19168 25740 19174
rect 25688 19110 25740 19116
rect 25594 18864 25650 18873
rect 25320 18828 25372 18834
rect 25594 18799 25650 18808
rect 25320 18770 25372 18776
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 24952 17128 25004 17134
rect 24952 17070 25004 17076
rect 24768 16516 24820 16522
rect 23020 16040 23072 16046
rect 23020 15982 23072 15988
rect 23480 16040 23532 16046
rect 23480 15982 23532 15988
rect 22744 15972 22796 15978
rect 22744 15914 22796 15920
rect 22468 15088 22520 15094
rect 22468 15030 22520 15036
rect 22480 14006 22508 15030
rect 22468 14000 22520 14006
rect 22468 13942 22520 13948
rect 22480 13258 22508 13942
rect 22756 13394 22784 15914
rect 23032 14550 23060 15982
rect 23097 15804 23393 15824
rect 23153 15802 23177 15804
rect 23233 15802 23257 15804
rect 23313 15802 23337 15804
rect 23175 15750 23177 15802
rect 23239 15750 23251 15802
rect 23313 15750 23315 15802
rect 23153 15748 23177 15750
rect 23233 15748 23257 15750
rect 23313 15748 23337 15750
rect 23097 15728 23393 15748
rect 23492 15706 23520 15982
rect 23480 15700 23532 15706
rect 23480 15642 23532 15648
rect 23097 14716 23393 14736
rect 23153 14714 23177 14716
rect 23233 14714 23257 14716
rect 23313 14714 23337 14716
rect 23175 14662 23177 14714
rect 23239 14662 23251 14714
rect 23313 14662 23315 14714
rect 23153 14660 23177 14662
rect 23233 14660 23257 14662
rect 23313 14660 23337 14662
rect 23097 14640 23393 14660
rect 23020 14544 23072 14550
rect 23020 14486 23072 14492
rect 23204 14340 23256 14346
rect 23204 14282 23256 14288
rect 23216 13802 23244 14282
rect 22928 13796 22980 13802
rect 22928 13738 22980 13744
rect 23204 13796 23256 13802
rect 23204 13738 23256 13744
rect 22836 13728 22888 13734
rect 22836 13670 22888 13676
rect 22848 13394 22876 13670
rect 22940 13530 22968 13738
rect 23097 13628 23393 13648
rect 23153 13626 23177 13628
rect 23233 13626 23257 13628
rect 23313 13626 23337 13628
rect 23175 13574 23177 13626
rect 23239 13574 23251 13626
rect 23313 13574 23315 13626
rect 23153 13572 23177 13574
rect 23233 13572 23257 13574
rect 23313 13572 23337 13574
rect 23097 13552 23393 13572
rect 22928 13524 22980 13530
rect 22928 13466 22980 13472
rect 22744 13388 22796 13394
rect 22744 13330 22796 13336
rect 22836 13388 22888 13394
rect 22836 13330 22888 13336
rect 22468 13252 22520 13258
rect 22468 13194 22520 13200
rect 22480 12918 22508 13194
rect 22468 12912 22520 12918
rect 22468 12854 22520 12860
rect 23572 12844 23624 12850
rect 23572 12786 23624 12792
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 23020 12776 23072 12782
rect 23020 12718 23072 12724
rect 22376 12708 22428 12714
rect 22376 12650 22428 12656
rect 22008 12368 22060 12374
rect 22008 12310 22060 12316
rect 22664 12238 22692 12718
rect 22744 12640 22796 12646
rect 22744 12582 22796 12588
rect 22756 12374 22784 12582
rect 23032 12442 23060 12718
rect 23097 12540 23393 12560
rect 23153 12538 23177 12540
rect 23233 12538 23257 12540
rect 23313 12538 23337 12540
rect 23175 12486 23177 12538
rect 23239 12486 23251 12538
rect 23313 12486 23315 12538
rect 23153 12484 23177 12486
rect 23233 12484 23257 12486
rect 23313 12484 23337 12486
rect 23097 12464 23393 12484
rect 23584 12442 23612 12786
rect 23020 12436 23072 12442
rect 23020 12378 23072 12384
rect 23572 12436 23624 12442
rect 23572 12378 23624 12384
rect 22744 12368 22796 12374
rect 22744 12310 22796 12316
rect 23112 12368 23164 12374
rect 23112 12310 23164 12316
rect 23124 12238 23152 12310
rect 22652 12232 22704 12238
rect 22652 12174 22704 12180
rect 23112 12232 23164 12238
rect 23112 12174 23164 12180
rect 23124 11642 23152 12174
rect 23032 11614 23152 11642
rect 23032 11354 23060 11614
rect 23572 11552 23624 11558
rect 23572 11494 23624 11500
rect 23097 11452 23393 11472
rect 23153 11450 23177 11452
rect 23233 11450 23257 11452
rect 23313 11450 23337 11452
rect 23175 11398 23177 11450
rect 23239 11398 23251 11450
rect 23313 11398 23315 11450
rect 23153 11396 23177 11398
rect 23233 11396 23257 11398
rect 23313 11396 23337 11398
rect 23097 11376 23393 11396
rect 23020 11348 23072 11354
rect 23020 11290 23072 11296
rect 23584 11218 23612 11494
rect 21732 11212 21784 11218
rect 21732 11154 21784 11160
rect 22376 11212 22428 11218
rect 22376 11154 22428 11160
rect 22560 11212 22612 11218
rect 22560 11154 22612 11160
rect 22836 11212 22888 11218
rect 22836 11154 22888 11160
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 21548 11076 21600 11082
rect 21548 11018 21600 11024
rect 21916 11076 21968 11082
rect 21916 11018 21968 11024
rect 21560 9518 21588 11018
rect 21928 9586 21956 11018
rect 22388 10062 22416 11154
rect 22572 10266 22600 11154
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 22376 10056 22428 10062
rect 22376 9998 22428 10004
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 21548 9512 21600 9518
rect 21548 9454 21600 9460
rect 22388 9178 22416 9998
rect 22572 9518 22600 10202
rect 22848 9926 22876 11154
rect 23480 11076 23532 11082
rect 23480 11018 23532 11024
rect 23020 10464 23072 10470
rect 23020 10406 23072 10412
rect 23032 10130 23060 10406
rect 23097 10364 23393 10384
rect 23153 10362 23177 10364
rect 23233 10362 23257 10364
rect 23313 10362 23337 10364
rect 23175 10310 23177 10362
rect 23239 10310 23251 10362
rect 23313 10310 23315 10362
rect 23153 10308 23177 10310
rect 23233 10308 23257 10310
rect 23313 10308 23337 10310
rect 23097 10288 23393 10308
rect 23020 10124 23072 10130
rect 23020 10066 23072 10072
rect 22836 9920 22888 9926
rect 22836 9862 22888 9868
rect 22560 9512 22612 9518
rect 22560 9454 22612 9460
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22100 8968 22152 8974
rect 22100 8910 22152 8916
rect 22112 8430 22140 8910
rect 22100 8424 22152 8430
rect 22100 8366 22152 8372
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 21652 7546 21680 7890
rect 22388 7834 22416 9114
rect 22848 8430 22876 9862
rect 23097 9276 23393 9296
rect 23153 9274 23177 9276
rect 23233 9274 23257 9276
rect 23313 9274 23337 9276
rect 23175 9222 23177 9274
rect 23239 9222 23251 9274
rect 23313 9222 23315 9274
rect 23153 9220 23177 9222
rect 23233 9220 23257 9222
rect 23313 9220 23337 9222
rect 23097 9200 23393 9220
rect 23492 8906 23520 11018
rect 23572 9444 23624 9450
rect 23572 9386 23624 9392
rect 23584 9178 23612 9386
rect 23572 9172 23624 9178
rect 23572 9114 23624 9120
rect 23572 8968 23624 8974
rect 23572 8910 23624 8916
rect 23480 8900 23532 8906
rect 23480 8842 23532 8848
rect 22836 8424 22888 8430
rect 22836 8366 22888 8372
rect 22560 8356 22612 8362
rect 22560 8298 22612 8304
rect 22928 8356 22980 8362
rect 22928 8298 22980 8304
rect 22296 7806 22416 7834
rect 21640 7540 21692 7546
rect 21640 7482 21692 7488
rect 22296 7342 22324 7806
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22388 7478 22416 7686
rect 22376 7472 22428 7478
rect 22376 7414 22428 7420
rect 21416 7296 21496 7324
rect 22284 7336 22336 7342
rect 21364 7278 21416 7284
rect 22284 7278 22336 7284
rect 22480 7274 22508 7686
rect 22468 7268 22520 7274
rect 22468 7210 22520 7216
rect 21272 6860 21324 6866
rect 21272 6802 21324 6808
rect 21732 6656 21784 6662
rect 21732 6598 21784 6604
rect 21744 6458 21772 6598
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 21732 6452 21784 6458
rect 21732 6394 21784 6400
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 21376 5778 21404 6054
rect 21364 5772 21416 5778
rect 21364 5714 21416 5720
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20628 4548 20680 4554
rect 20628 4490 20680 4496
rect 20732 4010 20760 4558
rect 20824 4282 20852 5170
rect 21376 5166 21404 5714
rect 21744 5642 21772 6394
rect 22480 6186 22508 7210
rect 22572 6730 22600 8298
rect 22940 7342 22968 8298
rect 23480 8288 23532 8294
rect 23480 8230 23532 8236
rect 23097 8188 23393 8208
rect 23153 8186 23177 8188
rect 23233 8186 23257 8188
rect 23313 8186 23337 8188
rect 23175 8134 23177 8186
rect 23239 8134 23251 8186
rect 23313 8134 23315 8186
rect 23153 8132 23177 8134
rect 23233 8132 23257 8134
rect 23313 8132 23337 8134
rect 23097 8112 23393 8132
rect 23492 7410 23520 8230
rect 23584 7546 23612 8910
rect 23572 7540 23624 7546
rect 23572 7482 23624 7488
rect 23480 7404 23532 7410
rect 23480 7346 23532 7352
rect 22928 7336 22980 7342
rect 22928 7278 22980 7284
rect 22928 7200 22980 7206
rect 22928 7142 22980 7148
rect 22560 6724 22612 6730
rect 22560 6666 22612 6672
rect 22572 6458 22600 6666
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 22468 6180 22520 6186
rect 22468 6122 22520 6128
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22572 5846 22600 6054
rect 22192 5840 22244 5846
rect 22192 5782 22244 5788
rect 22560 5840 22612 5846
rect 22560 5782 22612 5788
rect 21732 5636 21784 5642
rect 21732 5578 21784 5584
rect 22204 5370 22232 5782
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 22940 5166 22968 7142
rect 23097 7100 23393 7120
rect 23153 7098 23177 7100
rect 23233 7098 23257 7100
rect 23313 7098 23337 7100
rect 23175 7046 23177 7098
rect 23239 7046 23251 7098
rect 23313 7046 23315 7098
rect 23153 7044 23177 7046
rect 23233 7044 23257 7046
rect 23313 7044 23337 7046
rect 23097 7024 23393 7044
rect 23492 6866 23520 7346
rect 23480 6860 23532 6866
rect 23480 6802 23532 6808
rect 23676 6322 23704 16510
rect 24768 16458 24820 16464
rect 23940 15360 23992 15366
rect 23940 15302 23992 15308
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 23768 13326 23796 14214
rect 23756 13320 23808 13326
rect 23756 13262 23808 13268
rect 23848 11144 23900 11150
rect 23848 11086 23900 11092
rect 23756 11008 23808 11014
rect 23756 10950 23808 10956
rect 23768 10606 23796 10950
rect 23756 10600 23808 10606
rect 23756 10542 23808 10548
rect 23860 10266 23888 11086
rect 23848 10260 23900 10266
rect 23848 10202 23900 10208
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 23860 9042 23888 9318
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23848 8900 23900 8906
rect 23848 8842 23900 8848
rect 23756 8288 23808 8294
rect 23756 8230 23808 8236
rect 23768 7954 23796 8230
rect 23756 7948 23808 7954
rect 23756 7890 23808 7896
rect 23768 7342 23796 7890
rect 23860 7818 23888 8842
rect 23848 7812 23900 7818
rect 23848 7754 23900 7760
rect 23756 7336 23808 7342
rect 23756 7278 23808 7284
rect 23860 6798 23888 7754
rect 23952 6866 23980 15302
rect 24964 15162 24992 17070
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24400 14476 24452 14482
rect 24400 14418 24452 14424
rect 24412 13938 24440 14418
rect 24964 14278 24992 15098
rect 24952 14272 25004 14278
rect 24952 14214 25004 14220
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 24124 13320 24176 13326
rect 24124 13262 24176 13268
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 24044 12850 24072 13126
rect 24032 12844 24084 12850
rect 24032 12786 24084 12792
rect 24136 12442 24164 13262
rect 24124 12436 24176 12442
rect 24124 12378 24176 12384
rect 24412 9518 24440 13874
rect 25044 13796 25096 13802
rect 25044 13738 25096 13744
rect 25056 12986 25084 13738
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 25056 12714 25084 12922
rect 25044 12708 25096 12714
rect 25044 12650 25096 12656
rect 24860 12640 24912 12646
rect 24860 12582 24912 12588
rect 24872 12306 24900 12582
rect 24860 12300 24912 12306
rect 24860 12242 24912 12248
rect 24872 11694 24900 12242
rect 25056 11694 25084 12650
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 25044 11688 25096 11694
rect 25044 11630 25096 11636
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24596 9586 24624 10610
rect 24584 9580 24636 9586
rect 24584 9522 24636 9528
rect 24400 9512 24452 9518
rect 24400 9454 24452 9460
rect 24860 8356 24912 8362
rect 24860 8298 24912 8304
rect 24872 8090 24900 8298
rect 24860 8084 24912 8090
rect 24860 8026 24912 8032
rect 24124 7880 24176 7886
rect 24124 7822 24176 7828
rect 24136 7546 24164 7822
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 23940 6860 23992 6866
rect 23940 6802 23992 6808
rect 23848 6792 23900 6798
rect 23848 6734 23900 6740
rect 24032 6792 24084 6798
rect 24032 6734 24084 6740
rect 23020 6316 23072 6322
rect 23020 6258 23072 6264
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 23032 5370 23060 6258
rect 23097 6012 23393 6032
rect 23153 6010 23177 6012
rect 23233 6010 23257 6012
rect 23313 6010 23337 6012
rect 23175 5958 23177 6010
rect 23239 5958 23251 6010
rect 23313 5958 23315 6010
rect 23153 5956 23177 5958
rect 23233 5956 23257 5958
rect 23313 5956 23337 5958
rect 23097 5936 23393 5956
rect 23480 5568 23532 5574
rect 23480 5510 23532 5516
rect 23020 5364 23072 5370
rect 23020 5306 23072 5312
rect 23492 5166 23520 5510
rect 24044 5370 24072 6734
rect 24400 6656 24452 6662
rect 24400 6598 24452 6604
rect 24412 6254 24440 6598
rect 24400 6248 24452 6254
rect 24400 6190 24452 6196
rect 24308 5772 24360 5778
rect 24308 5714 24360 5720
rect 24032 5364 24084 5370
rect 24032 5306 24084 5312
rect 24320 5166 24348 5714
rect 21364 5160 21416 5166
rect 21364 5102 21416 5108
rect 22928 5160 22980 5166
rect 22928 5102 22980 5108
rect 23480 5160 23532 5166
rect 23480 5102 23532 5108
rect 24308 5160 24360 5166
rect 24308 5102 24360 5108
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20916 4758 20944 4966
rect 23097 4924 23393 4944
rect 23153 4922 23177 4924
rect 23233 4922 23257 4924
rect 23313 4922 23337 4924
rect 23175 4870 23177 4922
rect 23239 4870 23251 4922
rect 23313 4870 23315 4922
rect 23153 4868 23177 4870
rect 23233 4868 23257 4870
rect 23313 4868 23337 4870
rect 23097 4848 23393 4868
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 20904 4752 20956 4758
rect 20904 4694 20956 4700
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 20812 4276 20864 4282
rect 20812 4218 20864 4224
rect 21008 4078 21036 4422
rect 22388 4146 22416 4762
rect 24400 4684 24452 4690
rect 24400 4626 24452 4632
rect 22928 4480 22980 4486
rect 22928 4422 22980 4428
rect 22940 4282 22968 4422
rect 22928 4276 22980 4282
rect 22928 4218 22980 4224
rect 21088 4140 21140 4146
rect 21088 4082 21140 4088
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 20996 4072 21048 4078
rect 20996 4014 21048 4020
rect 20720 4004 20772 4010
rect 20720 3946 20772 3952
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 20456 2990 20484 3334
rect 20444 2984 20496 2990
rect 20732 2938 20760 3946
rect 21100 3602 21128 4082
rect 24412 3942 24440 4626
rect 24400 3936 24452 3942
rect 24400 3878 24452 3884
rect 23097 3836 23393 3856
rect 23153 3834 23177 3836
rect 23233 3834 23257 3836
rect 23313 3834 23337 3836
rect 23175 3782 23177 3834
rect 23239 3782 23251 3834
rect 23313 3782 23315 3834
rect 23153 3780 23177 3782
rect 23233 3780 23257 3782
rect 23313 3780 23337 3782
rect 23097 3760 23393 3780
rect 21088 3596 21140 3602
rect 21088 3538 21140 3544
rect 20444 2926 20496 2932
rect 19892 2916 19944 2922
rect 19892 2858 19944 2864
rect 20548 2910 20760 2938
rect 21916 2984 21968 2990
rect 21916 2926 21968 2932
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 17592 2644 17644 2650
rect 17592 2586 17644 2592
rect 18420 2644 18472 2650
rect 18420 2586 18472 2592
rect 19444 2582 19472 2790
rect 19904 2774 19932 2858
rect 20548 2854 20576 2910
rect 20536 2848 20588 2854
rect 20536 2790 20588 2796
rect 20720 2848 20772 2854
rect 20720 2790 20772 2796
rect 19904 2746 20024 2774
rect 16488 2576 16540 2582
rect 16488 2518 16540 2524
rect 19432 2576 19484 2582
rect 19432 2518 19484 2524
rect 19996 2446 20024 2746
rect 20548 2514 20576 2790
rect 20732 2582 20760 2790
rect 21928 2650 21956 2926
rect 25148 2774 25176 17274
rect 25228 16652 25280 16658
rect 25228 16594 25280 16600
rect 25240 16114 25268 16594
rect 25228 16108 25280 16114
rect 25228 16050 25280 16056
rect 25332 15978 25360 18770
rect 25412 18624 25464 18630
rect 25412 18566 25464 18572
rect 25424 18222 25452 18566
rect 25412 18216 25464 18222
rect 25412 18158 25464 18164
rect 25608 17202 25636 18799
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25700 16998 25728 19110
rect 25688 16992 25740 16998
rect 25688 16934 25740 16940
rect 25700 16658 25728 16934
rect 25688 16652 25740 16658
rect 25688 16594 25740 16600
rect 25596 16040 25648 16046
rect 25700 16028 25728 16594
rect 25648 16000 25728 16028
rect 25596 15982 25648 15988
rect 25320 15972 25372 15978
rect 25320 15914 25372 15920
rect 25700 15570 25728 16000
rect 25688 15564 25740 15570
rect 25688 15506 25740 15512
rect 25228 15496 25280 15502
rect 25228 15438 25280 15444
rect 25240 14618 25268 15438
rect 25320 15360 25372 15366
rect 25320 15302 25372 15308
rect 25332 14958 25360 15302
rect 25792 15162 25820 19858
rect 26068 18714 26096 20538
rect 26160 18834 26188 20946
rect 26436 20942 26464 21354
rect 26528 21010 26556 21830
rect 26516 21004 26568 21010
rect 26516 20946 26568 20952
rect 26424 20936 26476 20942
rect 26620 20890 26648 27950
rect 26712 27538 26740 31962
rect 27816 31278 27844 32302
rect 29196 32286 29316 32314
rect 29196 31754 29224 32286
rect 29276 32224 29328 32230
rect 29276 32166 29328 32172
rect 29288 31958 29316 32166
rect 29276 31952 29328 31958
rect 29276 31894 29328 31900
rect 29472 31822 29500 32370
rect 30024 31958 30052 33322
rect 30472 32292 30524 32298
rect 30472 32234 30524 32240
rect 30656 32292 30708 32298
rect 30656 32234 30708 32240
rect 30484 32026 30512 32234
rect 30472 32020 30524 32026
rect 30472 31962 30524 31968
rect 30012 31952 30064 31958
rect 30012 31894 30064 31900
rect 29552 31884 29604 31890
rect 29552 31826 29604 31832
rect 29460 31816 29512 31822
rect 29460 31758 29512 31764
rect 29196 31748 29420 31754
rect 29196 31726 29368 31748
rect 29368 31690 29420 31696
rect 28080 31680 28132 31686
rect 28080 31622 28132 31628
rect 28092 31346 28120 31622
rect 28632 31580 28928 31600
rect 28688 31578 28712 31580
rect 28768 31578 28792 31580
rect 28848 31578 28872 31580
rect 28710 31526 28712 31578
rect 28774 31526 28786 31578
rect 28848 31526 28850 31578
rect 28688 31524 28712 31526
rect 28768 31524 28792 31526
rect 28848 31524 28872 31526
rect 28632 31504 28928 31524
rect 28080 31340 28132 31346
rect 28080 31282 28132 31288
rect 27620 31272 27672 31278
rect 27620 31214 27672 31220
rect 27804 31272 27856 31278
rect 27804 31214 27856 31220
rect 27632 30802 27660 31214
rect 29380 31210 29408 31690
rect 29368 31204 29420 31210
rect 29368 31146 29420 31152
rect 27620 30796 27672 30802
rect 27620 30738 27672 30744
rect 27344 30728 27396 30734
rect 27344 30670 27396 30676
rect 27356 30326 27384 30670
rect 27344 30320 27396 30326
rect 27344 30262 27396 30268
rect 27632 29646 27660 30738
rect 28632 30492 28928 30512
rect 28688 30490 28712 30492
rect 28768 30490 28792 30492
rect 28848 30490 28872 30492
rect 28710 30438 28712 30490
rect 28774 30438 28786 30490
rect 28848 30438 28850 30490
rect 28688 30436 28712 30438
rect 28768 30436 28792 30438
rect 28848 30436 28872 30438
rect 28632 30416 28928 30436
rect 28356 30252 28408 30258
rect 28356 30194 28408 30200
rect 28368 29714 28396 30194
rect 28356 29708 28408 29714
rect 28356 29650 28408 29656
rect 29000 29708 29052 29714
rect 29000 29650 29052 29656
rect 27620 29640 27672 29646
rect 27620 29582 27672 29588
rect 27632 29238 27660 29582
rect 27896 29572 27948 29578
rect 27896 29514 27948 29520
rect 27620 29232 27672 29238
rect 27620 29174 27672 29180
rect 27632 28626 27660 29174
rect 27620 28620 27672 28626
rect 27620 28562 27672 28568
rect 27632 28082 27660 28562
rect 27620 28076 27672 28082
rect 27620 28018 27672 28024
rect 26700 27532 26752 27538
rect 26700 27474 26752 27480
rect 27632 27062 27660 28018
rect 27620 27056 27672 27062
rect 27620 26998 27672 27004
rect 27632 26382 27660 26998
rect 27804 26920 27856 26926
rect 27804 26862 27856 26868
rect 27816 26586 27844 26862
rect 27804 26580 27856 26586
rect 27804 26522 27856 26528
rect 27620 26376 27672 26382
rect 27620 26318 27672 26324
rect 27528 26036 27580 26042
rect 27528 25978 27580 25984
rect 26976 25832 27028 25838
rect 26896 25780 26976 25786
rect 26896 25774 27028 25780
rect 26896 25758 27016 25774
rect 26896 25294 26924 25758
rect 26884 25288 26936 25294
rect 26884 25230 26936 25236
rect 26896 24206 26924 25230
rect 27160 24608 27212 24614
rect 27160 24550 27212 24556
rect 27172 24342 27200 24550
rect 27160 24336 27212 24342
rect 27160 24278 27212 24284
rect 26884 24200 26936 24206
rect 26884 24142 26936 24148
rect 26896 23866 26924 24142
rect 26884 23860 26936 23866
rect 26884 23802 26936 23808
rect 26792 23520 26844 23526
rect 26792 23462 26844 23468
rect 26804 23254 26832 23462
rect 26792 23248 26844 23254
rect 26792 23190 26844 23196
rect 26424 20878 26476 20884
rect 26528 20862 26648 20890
rect 26424 20392 26476 20398
rect 26424 20334 26476 20340
rect 26436 19922 26464 20334
rect 26528 20058 26556 20862
rect 26608 20800 26660 20806
rect 26608 20742 26660 20748
rect 26620 20398 26648 20742
rect 26608 20392 26660 20398
rect 26608 20334 26660 20340
rect 26516 20052 26568 20058
rect 26516 19994 26568 20000
rect 26424 19916 26476 19922
rect 26424 19858 26476 19864
rect 26240 19168 26292 19174
rect 26240 19110 26292 19116
rect 26148 18828 26200 18834
rect 26148 18770 26200 18776
rect 25976 18698 26096 18714
rect 25964 18692 26096 18698
rect 26016 18686 26096 18692
rect 25964 18634 26016 18640
rect 25964 17060 26016 17066
rect 25964 17002 26016 17008
rect 25872 15632 25924 15638
rect 25872 15574 25924 15580
rect 25884 15162 25912 15574
rect 25780 15156 25832 15162
rect 25780 15098 25832 15104
rect 25872 15156 25924 15162
rect 25872 15098 25924 15104
rect 25320 14952 25372 14958
rect 25320 14894 25372 14900
rect 25228 14612 25280 14618
rect 25228 14554 25280 14560
rect 25792 14482 25820 15098
rect 25780 14476 25832 14482
rect 25780 14418 25832 14424
rect 25884 14346 25912 15098
rect 25872 14340 25924 14346
rect 25872 14282 25924 14288
rect 25596 14068 25648 14074
rect 25596 14010 25648 14016
rect 25608 12434 25636 14010
rect 25976 13734 26004 17002
rect 26068 16522 26096 18686
rect 26160 18426 26188 18770
rect 26148 18420 26200 18426
rect 26148 18362 26200 18368
rect 26252 17134 26280 19110
rect 26528 18970 26556 19994
rect 26620 19310 26648 20334
rect 26608 19304 26660 19310
rect 26608 19246 26660 19252
rect 26516 18964 26568 18970
rect 26516 18906 26568 18912
rect 26332 18896 26384 18902
rect 26332 18838 26384 18844
rect 26240 17128 26292 17134
rect 26240 17070 26292 17076
rect 26148 16992 26200 16998
rect 26148 16934 26200 16940
rect 26056 16516 26108 16522
rect 26056 16458 26108 16464
rect 26068 15638 26096 16458
rect 26056 15632 26108 15638
rect 26056 15574 26108 15580
rect 26056 15360 26108 15366
rect 26056 15302 26108 15308
rect 25964 13728 26016 13734
rect 25964 13670 26016 13676
rect 25976 12782 26004 13670
rect 26068 12986 26096 15302
rect 26160 14550 26188 16934
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 26252 16250 26280 16594
rect 26240 16244 26292 16250
rect 26240 16186 26292 16192
rect 26344 16046 26372 18838
rect 26424 17672 26476 17678
rect 26424 17614 26476 17620
rect 26436 16590 26464 17614
rect 26528 16794 26556 18906
rect 26700 18828 26752 18834
rect 26700 18770 26752 18776
rect 26712 17134 26740 18770
rect 26804 17814 26832 23190
rect 26896 22574 26924 23802
rect 27540 22982 27568 25978
rect 27908 24410 27936 29514
rect 28632 29404 28928 29424
rect 28688 29402 28712 29404
rect 28768 29402 28792 29404
rect 28848 29402 28872 29404
rect 28710 29350 28712 29402
rect 28774 29350 28786 29402
rect 28848 29350 28850 29402
rect 28688 29348 28712 29350
rect 28768 29348 28792 29350
rect 28848 29348 28872 29350
rect 28632 29328 28928 29348
rect 28264 29028 28316 29034
rect 28264 28970 28316 28976
rect 28276 28762 28304 28970
rect 29012 28762 29040 29650
rect 29380 29102 29408 31146
rect 29564 31142 29592 31826
rect 29920 31816 29972 31822
rect 29920 31758 29972 31764
rect 29552 31136 29604 31142
rect 29552 31078 29604 31084
rect 29564 30190 29592 31078
rect 29932 30258 29960 31758
rect 29920 30252 29972 30258
rect 29920 30194 29972 30200
rect 30024 30190 30052 31894
rect 30668 31754 30696 32234
rect 30748 32224 30800 32230
rect 30748 32166 30800 32172
rect 30760 32026 30788 32166
rect 30748 32020 30800 32026
rect 30748 31962 30800 31968
rect 31208 31816 31260 31822
rect 31208 31758 31260 31764
rect 31668 31816 31720 31822
rect 31668 31758 31720 31764
rect 30656 31748 30708 31754
rect 30656 31690 30708 31696
rect 30668 30938 30696 31690
rect 31220 31328 31248 31758
rect 31300 31340 31352 31346
rect 31220 31300 31300 31328
rect 31024 31136 31076 31142
rect 31024 31078 31076 31084
rect 30656 30932 30708 30938
rect 30656 30874 30708 30880
rect 31036 30870 31064 31078
rect 31024 30864 31076 30870
rect 31024 30806 31076 30812
rect 29552 30184 29604 30190
rect 29552 30126 29604 30132
rect 30012 30184 30064 30190
rect 30012 30126 30064 30132
rect 30932 29640 30984 29646
rect 30932 29582 30984 29588
rect 30944 29306 30972 29582
rect 30932 29300 30984 29306
rect 30932 29242 30984 29248
rect 31220 29170 31248 31300
rect 31300 31282 31352 31288
rect 31680 31278 31708 31758
rect 31668 31272 31720 31278
rect 31668 31214 31720 31220
rect 31300 31136 31352 31142
rect 31300 31078 31352 31084
rect 31312 29510 31340 31078
rect 31680 30938 31708 31214
rect 31668 30932 31720 30938
rect 31668 30874 31720 30880
rect 31484 30864 31536 30870
rect 31484 30806 31536 30812
rect 31496 30410 31524 30806
rect 31496 30382 31800 30410
rect 31772 29850 31800 30382
rect 31760 29844 31812 29850
rect 31760 29786 31812 29792
rect 31300 29504 31352 29510
rect 31300 29446 31352 29452
rect 31208 29164 31260 29170
rect 31208 29106 31260 29112
rect 29368 29096 29420 29102
rect 29368 29038 29420 29044
rect 30104 29096 30156 29102
rect 30104 29038 30156 29044
rect 28264 28756 28316 28762
rect 28264 28698 28316 28704
rect 29000 28756 29052 28762
rect 29000 28698 29052 28704
rect 29276 28552 29328 28558
rect 29276 28494 29328 28500
rect 28632 28316 28928 28336
rect 28688 28314 28712 28316
rect 28768 28314 28792 28316
rect 28848 28314 28872 28316
rect 28710 28262 28712 28314
rect 28774 28262 28786 28314
rect 28848 28262 28850 28314
rect 28688 28260 28712 28262
rect 28768 28260 28792 28262
rect 28848 28260 28872 28262
rect 28632 28240 28928 28260
rect 29288 28218 29316 28494
rect 29276 28212 29328 28218
rect 29276 28154 29328 28160
rect 30116 27946 30144 29038
rect 30288 29028 30340 29034
rect 30288 28970 30340 28976
rect 30300 28694 30328 28970
rect 30288 28688 30340 28694
rect 30288 28630 30340 28636
rect 30300 28558 30328 28630
rect 30288 28552 30340 28558
rect 30288 28494 30340 28500
rect 31220 28490 31248 29106
rect 31312 29102 31340 29446
rect 31300 29096 31352 29102
rect 31300 29038 31352 29044
rect 31312 28558 31340 29038
rect 31300 28552 31352 28558
rect 31300 28494 31352 28500
rect 31944 28552 31996 28558
rect 31944 28494 31996 28500
rect 31208 28484 31260 28490
rect 31208 28426 31260 28432
rect 31220 28218 31248 28426
rect 31208 28212 31260 28218
rect 31208 28154 31260 28160
rect 28724 27940 28776 27946
rect 28724 27882 28776 27888
rect 30104 27940 30156 27946
rect 30104 27882 30156 27888
rect 30380 27940 30432 27946
rect 30380 27882 30432 27888
rect 28736 27674 28764 27882
rect 28724 27668 28776 27674
rect 28724 27610 28776 27616
rect 28264 27532 28316 27538
rect 28264 27474 28316 27480
rect 28172 26784 28224 26790
rect 28172 26726 28224 26732
rect 28184 25362 28212 26726
rect 28172 25356 28224 25362
rect 28172 25298 28224 25304
rect 28184 24750 28212 25298
rect 28172 24744 28224 24750
rect 28172 24686 28224 24692
rect 28276 24614 28304 27474
rect 28632 27228 28928 27248
rect 28688 27226 28712 27228
rect 28768 27226 28792 27228
rect 28848 27226 28872 27228
rect 28710 27174 28712 27226
rect 28774 27174 28786 27226
rect 28848 27174 28850 27226
rect 28688 27172 28712 27174
rect 28768 27172 28792 27174
rect 28848 27172 28872 27174
rect 28632 27152 28928 27172
rect 29828 26988 29880 26994
rect 29828 26930 29880 26936
rect 29368 26240 29420 26246
rect 29368 26182 29420 26188
rect 28632 26140 28928 26160
rect 28688 26138 28712 26140
rect 28768 26138 28792 26140
rect 28848 26138 28872 26140
rect 28710 26086 28712 26138
rect 28774 26086 28786 26138
rect 28848 26086 28850 26138
rect 28688 26084 28712 26086
rect 28768 26084 28792 26086
rect 28848 26084 28872 26086
rect 28632 26064 28928 26084
rect 28448 25900 28500 25906
rect 28448 25842 28500 25848
rect 28460 25362 28488 25842
rect 28540 25764 28592 25770
rect 28540 25706 28592 25712
rect 28552 25498 28580 25706
rect 28540 25492 28592 25498
rect 28540 25434 28592 25440
rect 29380 25362 29408 26182
rect 29840 25770 29868 26930
rect 30116 26926 30144 27882
rect 30104 26920 30156 26926
rect 30104 26862 30156 26868
rect 30116 26518 30144 26862
rect 30104 26512 30156 26518
rect 30104 26454 30156 26460
rect 30392 26042 30420 27882
rect 30656 27872 30708 27878
rect 30656 27814 30708 27820
rect 30668 27538 30696 27814
rect 30656 27532 30708 27538
rect 30656 27474 30708 27480
rect 31956 27470 31984 28494
rect 31944 27464 31996 27470
rect 31772 27412 31944 27418
rect 31772 27406 31996 27412
rect 30472 27396 30524 27402
rect 30472 27338 30524 27344
rect 31772 27390 31984 27406
rect 30380 26036 30432 26042
rect 30380 25978 30432 25984
rect 29828 25764 29880 25770
rect 29828 25706 29880 25712
rect 28448 25356 28500 25362
rect 28448 25298 28500 25304
rect 29368 25356 29420 25362
rect 29368 25298 29420 25304
rect 28264 24608 28316 24614
rect 28264 24550 28316 24556
rect 28356 24608 28408 24614
rect 28356 24550 28408 24556
rect 27896 24404 27948 24410
rect 27896 24346 27948 24352
rect 28172 23520 28224 23526
rect 28172 23462 28224 23468
rect 28184 23186 28212 23462
rect 28276 23254 28304 24550
rect 28368 24206 28396 24550
rect 28460 24342 28488 25298
rect 28632 25052 28928 25072
rect 28688 25050 28712 25052
rect 28768 25050 28792 25052
rect 28848 25050 28872 25052
rect 28710 24998 28712 25050
rect 28774 24998 28786 25050
rect 28848 24998 28850 25050
rect 28688 24996 28712 24998
rect 28768 24996 28792 24998
rect 28848 24996 28872 24998
rect 28632 24976 28928 24996
rect 29184 24744 29236 24750
rect 29184 24686 29236 24692
rect 29196 24410 29224 24686
rect 29184 24404 29236 24410
rect 29184 24346 29236 24352
rect 28448 24336 28500 24342
rect 28448 24278 28500 24284
rect 28356 24200 28408 24206
rect 28356 24142 28408 24148
rect 28460 23730 28488 24278
rect 28540 24200 28592 24206
rect 28540 24142 28592 24148
rect 28448 23724 28500 23730
rect 28448 23666 28500 23672
rect 28552 23662 28580 24142
rect 29840 24138 29868 25706
rect 30484 24970 30512 27338
rect 30564 27328 30616 27334
rect 30564 27270 30616 27276
rect 31208 27328 31260 27334
rect 31208 27270 31260 27276
rect 30576 26382 30604 27270
rect 30564 26376 30616 26382
rect 30564 26318 30616 26324
rect 30932 25968 30984 25974
rect 30932 25910 30984 25916
rect 30748 25832 30800 25838
rect 30748 25774 30800 25780
rect 30484 24942 30604 24970
rect 30760 24954 30788 25774
rect 30472 24812 30524 24818
rect 30472 24754 30524 24760
rect 29828 24132 29880 24138
rect 29828 24074 29880 24080
rect 28632 23964 28928 23984
rect 28688 23962 28712 23964
rect 28768 23962 28792 23964
rect 28848 23962 28872 23964
rect 28710 23910 28712 23962
rect 28774 23910 28786 23962
rect 28848 23910 28850 23962
rect 28688 23908 28712 23910
rect 28768 23908 28792 23910
rect 28848 23908 28872 23910
rect 28632 23888 28928 23908
rect 29460 23792 29512 23798
rect 29460 23734 29512 23740
rect 28540 23656 28592 23662
rect 28540 23598 28592 23604
rect 28448 23316 28500 23322
rect 28448 23258 28500 23264
rect 28264 23248 28316 23254
rect 28264 23190 28316 23196
rect 28172 23180 28224 23186
rect 28172 23122 28224 23128
rect 27804 23044 27856 23050
rect 27804 22986 27856 22992
rect 27528 22976 27580 22982
rect 27528 22918 27580 22924
rect 27540 22642 27568 22918
rect 27068 22636 27120 22642
rect 27068 22578 27120 22584
rect 27528 22636 27580 22642
rect 27528 22578 27580 22584
rect 26884 22568 26936 22574
rect 26884 22510 26936 22516
rect 27080 22098 27108 22578
rect 27068 22092 27120 22098
rect 27068 22034 27120 22040
rect 27436 22092 27488 22098
rect 27436 22034 27488 22040
rect 27080 21554 27108 22034
rect 27252 21616 27304 21622
rect 27252 21558 27304 21564
rect 27068 21548 27120 21554
rect 27068 21490 27120 21496
rect 27264 21010 27292 21558
rect 27448 21078 27476 22034
rect 27436 21072 27488 21078
rect 27436 21014 27488 21020
rect 27252 21004 27304 21010
rect 27252 20946 27304 20952
rect 27264 20534 27292 20946
rect 27620 20800 27672 20806
rect 27620 20742 27672 20748
rect 27252 20528 27304 20534
rect 27252 20470 27304 20476
rect 27632 20262 27660 20742
rect 27620 20256 27672 20262
rect 27620 20198 27672 20204
rect 27632 19990 27660 20198
rect 27620 19984 27672 19990
rect 27620 19926 27672 19932
rect 27252 19916 27304 19922
rect 27252 19858 27304 19864
rect 27344 19916 27396 19922
rect 27344 19858 27396 19864
rect 27264 19514 27292 19858
rect 27252 19508 27304 19514
rect 27252 19450 27304 19456
rect 26976 19236 27028 19242
rect 26976 19178 27028 19184
rect 26792 17808 26844 17814
rect 26792 17750 26844 17756
rect 26700 17128 26752 17134
rect 26700 17070 26752 17076
rect 26516 16788 26568 16794
rect 26568 16748 26648 16776
rect 26516 16730 26568 16736
rect 26424 16584 26476 16590
rect 26424 16526 26476 16532
rect 26516 16448 26568 16454
rect 26516 16390 26568 16396
rect 26332 16040 26384 16046
rect 26332 15982 26384 15988
rect 26344 15502 26372 15982
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 26528 14958 26556 16390
rect 26620 15570 26648 16748
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26516 14952 26568 14958
rect 26516 14894 26568 14900
rect 26620 14618 26648 15506
rect 26792 15360 26844 15366
rect 26792 15302 26844 15308
rect 26804 15026 26832 15302
rect 26792 15020 26844 15026
rect 26792 14962 26844 14968
rect 26608 14612 26660 14618
rect 26528 14572 26608 14600
rect 26148 14544 26200 14550
rect 26148 14486 26200 14492
rect 26160 13394 26188 14486
rect 26528 13870 26556 14572
rect 26608 14554 26660 14560
rect 26608 14408 26660 14414
rect 26608 14350 26660 14356
rect 26620 14074 26648 14350
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26516 13864 26568 13870
rect 26516 13806 26568 13812
rect 26988 13462 27016 19178
rect 27264 18834 27292 19450
rect 27356 19310 27384 19858
rect 27344 19304 27396 19310
rect 27344 19246 27396 19252
rect 27252 18828 27304 18834
rect 27252 18770 27304 18776
rect 27160 18624 27212 18630
rect 27160 18566 27212 18572
rect 27172 18290 27200 18566
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 27632 17814 27660 19926
rect 27816 18426 27844 22986
rect 28184 22166 28212 23122
rect 28276 22778 28304 23190
rect 28264 22772 28316 22778
rect 28264 22714 28316 22720
rect 28172 22160 28224 22166
rect 28172 22102 28224 22108
rect 27988 22024 28040 22030
rect 27988 21966 28040 21972
rect 28000 21486 28028 21966
rect 28184 21486 28212 22102
rect 27988 21480 28040 21486
rect 27988 21422 28040 21428
rect 28172 21480 28224 21486
rect 28172 21422 28224 21428
rect 28264 20460 28316 20466
rect 28264 20402 28316 20408
rect 28276 19854 28304 20402
rect 28460 20398 28488 23258
rect 29368 23180 29420 23186
rect 29368 23122 29420 23128
rect 28540 22976 28592 22982
rect 28540 22918 28592 22924
rect 28552 22642 28580 22918
rect 28632 22876 28928 22896
rect 28688 22874 28712 22876
rect 28768 22874 28792 22876
rect 28848 22874 28872 22876
rect 28710 22822 28712 22874
rect 28774 22822 28786 22874
rect 28848 22822 28850 22874
rect 28688 22820 28712 22822
rect 28768 22820 28792 22822
rect 28848 22820 28872 22822
rect 28632 22800 28928 22820
rect 28540 22636 28592 22642
rect 28540 22578 28592 22584
rect 29380 22438 29408 23122
rect 29368 22432 29420 22438
rect 29368 22374 29420 22380
rect 28632 21788 28928 21808
rect 28688 21786 28712 21788
rect 28768 21786 28792 21788
rect 28848 21786 28872 21788
rect 28710 21734 28712 21786
rect 28774 21734 28786 21786
rect 28848 21734 28850 21786
rect 28688 21732 28712 21734
rect 28768 21732 28792 21734
rect 28848 21732 28872 21734
rect 28632 21712 28928 21732
rect 29000 21344 29052 21350
rect 29000 21286 29052 21292
rect 28632 20700 28928 20720
rect 28688 20698 28712 20700
rect 28768 20698 28792 20700
rect 28848 20698 28872 20700
rect 28710 20646 28712 20698
rect 28774 20646 28786 20698
rect 28848 20646 28850 20698
rect 28688 20644 28712 20646
rect 28768 20644 28792 20646
rect 28848 20644 28872 20646
rect 28632 20624 28928 20644
rect 29012 20466 29040 21286
rect 29092 21004 29144 21010
rect 29092 20946 29144 20952
rect 29104 20602 29132 20946
rect 29380 20942 29408 22374
rect 29472 21690 29500 23734
rect 29644 23656 29696 23662
rect 29644 23598 29696 23604
rect 29656 21894 29684 23598
rect 29840 22778 29868 24074
rect 30484 23662 30512 24754
rect 30472 23656 30524 23662
rect 30472 23598 30524 23604
rect 30012 23044 30064 23050
rect 30012 22986 30064 22992
rect 30024 22778 30052 22986
rect 29828 22772 29880 22778
rect 29828 22714 29880 22720
rect 30012 22772 30064 22778
rect 30012 22714 30064 22720
rect 29840 22506 29868 22714
rect 29828 22500 29880 22506
rect 29828 22442 29880 22448
rect 29644 21888 29696 21894
rect 29644 21830 29696 21836
rect 29460 21684 29512 21690
rect 29460 21626 29512 21632
rect 29368 20936 29420 20942
rect 29368 20878 29420 20884
rect 29828 20936 29880 20942
rect 29828 20878 29880 20884
rect 29092 20596 29144 20602
rect 29092 20538 29144 20544
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 28448 20392 28500 20398
rect 28448 20334 28500 20340
rect 29840 20330 29868 20878
rect 30472 20800 30524 20806
rect 30472 20742 30524 20748
rect 30484 20466 30512 20742
rect 30472 20460 30524 20466
rect 30472 20402 30524 20408
rect 29828 20324 29880 20330
rect 29828 20266 29880 20272
rect 28264 19848 28316 19854
rect 28264 19790 28316 19796
rect 28448 19848 28500 19854
rect 28448 19790 28500 19796
rect 28460 19174 28488 19790
rect 29552 19712 29604 19718
rect 29552 19654 29604 19660
rect 28632 19612 28928 19632
rect 28688 19610 28712 19612
rect 28768 19610 28792 19612
rect 28848 19610 28872 19612
rect 28710 19558 28712 19610
rect 28774 19558 28786 19610
rect 28848 19558 28850 19610
rect 28688 19556 28712 19558
rect 28768 19556 28792 19558
rect 28848 19556 28872 19558
rect 28632 19536 28928 19556
rect 29564 19310 29592 19654
rect 29840 19310 29868 20266
rect 29552 19304 29604 19310
rect 29552 19246 29604 19252
rect 29828 19304 29880 19310
rect 29828 19246 29880 19252
rect 28448 19168 28500 19174
rect 28448 19110 28500 19116
rect 28460 18834 28488 19110
rect 29840 18834 29868 19246
rect 28172 18828 28224 18834
rect 28172 18770 28224 18776
rect 28448 18828 28500 18834
rect 28448 18770 28500 18776
rect 29828 18828 29880 18834
rect 29828 18770 29880 18776
rect 27896 18692 27948 18698
rect 27896 18634 27948 18640
rect 27804 18420 27856 18426
rect 27804 18362 27856 18368
rect 27804 18216 27856 18222
rect 27804 18158 27856 18164
rect 27620 17808 27672 17814
rect 27620 17750 27672 17756
rect 27816 17678 27844 18158
rect 27908 17882 27936 18634
rect 28080 18624 28132 18630
rect 28080 18566 28132 18572
rect 28092 18222 28120 18566
rect 28080 18216 28132 18222
rect 28080 18158 28132 18164
rect 27896 17876 27948 17882
rect 27896 17818 27948 17824
rect 27988 17740 28040 17746
rect 27988 17682 28040 17688
rect 27804 17672 27856 17678
rect 27804 17614 27856 17620
rect 28000 17134 28028 17682
rect 28184 17338 28212 18770
rect 28632 18524 28928 18544
rect 28688 18522 28712 18524
rect 28768 18522 28792 18524
rect 28848 18522 28872 18524
rect 28710 18470 28712 18522
rect 28774 18470 28786 18522
rect 28848 18470 28850 18522
rect 28688 18468 28712 18470
rect 28768 18468 28792 18470
rect 28848 18468 28872 18470
rect 28632 18448 28928 18468
rect 29840 18154 29868 18770
rect 30576 18426 30604 24942
rect 30748 24948 30800 24954
rect 30748 24890 30800 24896
rect 30760 24834 30788 24890
rect 30760 24806 30880 24834
rect 30944 24818 30972 25910
rect 30748 24744 30800 24750
rect 30748 24686 30800 24692
rect 30760 24070 30788 24686
rect 30852 24274 30880 24806
rect 30932 24812 30984 24818
rect 30932 24754 30984 24760
rect 31220 24410 31248 27270
rect 31772 27130 31800 27390
rect 31760 27124 31812 27130
rect 31760 27066 31812 27072
rect 31576 26852 31628 26858
rect 31576 26794 31628 26800
rect 31300 26444 31352 26450
rect 31300 26386 31352 26392
rect 31312 25838 31340 26386
rect 31300 25832 31352 25838
rect 31300 25774 31352 25780
rect 31392 25832 31444 25838
rect 31392 25774 31444 25780
rect 31404 25498 31432 25774
rect 31392 25492 31444 25498
rect 31392 25434 31444 25440
rect 31208 24404 31260 24410
rect 31208 24346 31260 24352
rect 30840 24268 30892 24274
rect 30840 24210 30892 24216
rect 31404 24206 31432 25434
rect 31588 25362 31616 26794
rect 31772 26382 31800 27066
rect 31760 26376 31812 26382
rect 31760 26318 31812 26324
rect 31760 26240 31812 26246
rect 31760 26182 31812 26188
rect 31668 25696 31720 25702
rect 31668 25638 31720 25644
rect 31680 25430 31708 25638
rect 31668 25424 31720 25430
rect 31668 25366 31720 25372
rect 31772 25362 31800 26182
rect 31576 25356 31628 25362
rect 31576 25298 31628 25304
rect 31760 25356 31812 25362
rect 31760 25298 31812 25304
rect 31852 25220 31904 25226
rect 31852 25162 31904 25168
rect 31864 24698 31892 25162
rect 31772 24682 31892 24698
rect 32128 24744 32180 24750
rect 32128 24686 32180 24692
rect 31760 24676 31892 24682
rect 31812 24670 31892 24676
rect 31760 24618 31812 24624
rect 31392 24200 31444 24206
rect 31392 24142 31444 24148
rect 31760 24200 31812 24206
rect 31760 24142 31812 24148
rect 30748 24064 30800 24070
rect 30748 24006 30800 24012
rect 30760 23730 30788 24006
rect 30748 23724 30800 23730
rect 30748 23666 30800 23672
rect 30656 23588 30708 23594
rect 30656 23530 30708 23536
rect 30668 21962 30696 23530
rect 31772 23322 31800 24142
rect 31864 23662 31892 24670
rect 32140 24342 32168 24686
rect 32128 24336 32180 24342
rect 32128 24278 32180 24284
rect 31852 23656 31904 23662
rect 31852 23598 31904 23604
rect 31760 23316 31812 23322
rect 31760 23258 31812 23264
rect 30932 23112 30984 23118
rect 30932 23054 30984 23060
rect 31024 23112 31076 23118
rect 31024 23054 31076 23060
rect 30944 22778 30972 23054
rect 30932 22772 30984 22778
rect 30932 22714 30984 22720
rect 31036 22658 31064 23054
rect 31392 22976 31444 22982
rect 31392 22918 31444 22924
rect 30840 22636 30892 22642
rect 30840 22578 30892 22584
rect 30944 22630 31064 22658
rect 31404 22642 31432 22918
rect 31392 22636 31444 22642
rect 30852 22166 30880 22578
rect 30944 22438 30972 22630
rect 31392 22578 31444 22584
rect 30932 22432 30984 22438
rect 30932 22374 30984 22380
rect 30840 22160 30892 22166
rect 30840 22102 30892 22108
rect 30656 21956 30708 21962
rect 30656 21898 30708 21904
rect 30564 18420 30616 18426
rect 30564 18362 30616 18368
rect 30668 18222 30696 21898
rect 30944 21894 30972 22374
rect 30932 21888 30984 21894
rect 30932 21830 30984 21836
rect 31404 21554 31432 22578
rect 31852 22160 31904 22166
rect 31852 22102 31904 22108
rect 31864 21554 31892 22102
rect 32036 22092 32088 22098
rect 32036 22034 32088 22040
rect 31208 21548 31260 21554
rect 31208 21490 31260 21496
rect 31392 21548 31444 21554
rect 31392 21490 31444 21496
rect 31852 21548 31904 21554
rect 31852 21490 31904 21496
rect 30840 21004 30892 21010
rect 30840 20946 30892 20952
rect 30852 20602 30880 20946
rect 31220 20942 31248 21490
rect 31208 20936 31260 20942
rect 31208 20878 31260 20884
rect 31760 20936 31812 20942
rect 31760 20878 31812 20884
rect 30840 20596 30892 20602
rect 30840 20538 30892 20544
rect 30852 19378 30880 20538
rect 31220 19378 31248 20878
rect 31772 19854 31800 20878
rect 32048 20602 32076 22034
rect 32220 21412 32272 21418
rect 32220 21354 32272 21360
rect 32128 21344 32180 21350
rect 32128 21286 32180 21292
rect 32140 21078 32168 21286
rect 32128 21072 32180 21078
rect 32128 21014 32180 21020
rect 32232 20942 32260 21354
rect 32220 20936 32272 20942
rect 32220 20878 32272 20884
rect 32036 20596 32088 20602
rect 32036 20538 32088 20544
rect 32232 20398 32260 20878
rect 32220 20392 32272 20398
rect 32220 20334 32272 20340
rect 31760 19848 31812 19854
rect 31760 19790 31812 19796
rect 32128 19848 32180 19854
rect 32128 19790 32180 19796
rect 30840 19372 30892 19378
rect 30840 19314 30892 19320
rect 31208 19372 31260 19378
rect 31208 19314 31260 19320
rect 30748 19168 30800 19174
rect 30748 19110 30800 19116
rect 30760 18902 30788 19110
rect 30748 18896 30800 18902
rect 30748 18838 30800 18844
rect 31220 18766 31248 19314
rect 31772 19310 31800 19790
rect 31760 19304 31812 19310
rect 31760 19246 31812 19252
rect 31208 18760 31260 18766
rect 31208 18702 31260 18708
rect 31576 18420 31628 18426
rect 31576 18362 31628 18368
rect 30656 18216 30708 18222
rect 30656 18158 30708 18164
rect 30932 18216 30984 18222
rect 30932 18158 30984 18164
rect 29828 18148 29880 18154
rect 29828 18090 29880 18096
rect 28264 17672 28316 17678
rect 28264 17614 28316 17620
rect 28172 17332 28224 17338
rect 28172 17274 28224 17280
rect 28276 17134 28304 17614
rect 28632 17436 28928 17456
rect 28688 17434 28712 17436
rect 28768 17434 28792 17436
rect 28848 17434 28872 17436
rect 28710 17382 28712 17434
rect 28774 17382 28786 17434
rect 28848 17382 28850 17434
rect 28688 17380 28712 17382
rect 28768 17380 28792 17382
rect 28848 17380 28872 17382
rect 28632 17360 28928 17380
rect 30288 17264 30340 17270
rect 30288 17206 30340 17212
rect 27988 17128 28040 17134
rect 27988 17070 28040 17076
rect 28264 17128 28316 17134
rect 28264 17070 28316 17076
rect 28000 15638 28028 17070
rect 28276 16250 28304 17070
rect 29092 17060 29144 17066
rect 29092 17002 29144 17008
rect 29000 16992 29052 16998
rect 29000 16934 29052 16940
rect 28540 16720 28592 16726
rect 28540 16662 28592 16668
rect 28264 16244 28316 16250
rect 28264 16186 28316 16192
rect 28552 16046 28580 16662
rect 28632 16348 28928 16368
rect 28688 16346 28712 16348
rect 28768 16346 28792 16348
rect 28848 16346 28872 16348
rect 28710 16294 28712 16346
rect 28774 16294 28786 16346
rect 28848 16294 28850 16346
rect 28688 16292 28712 16294
rect 28768 16292 28792 16294
rect 28848 16292 28872 16294
rect 28632 16272 28928 16292
rect 28540 16040 28592 16046
rect 28540 15982 28592 15988
rect 29012 16028 29040 16934
rect 29104 16250 29132 17002
rect 29092 16244 29144 16250
rect 29092 16186 29144 16192
rect 29184 16040 29236 16046
rect 29012 16000 29184 16028
rect 27988 15632 28040 15638
rect 27988 15574 28040 15580
rect 27712 15564 27764 15570
rect 27712 15506 27764 15512
rect 27620 15496 27672 15502
rect 27620 15438 27672 15444
rect 27632 15026 27660 15438
rect 27724 15162 27752 15506
rect 27712 15156 27764 15162
rect 27712 15098 27764 15104
rect 27620 15020 27672 15026
rect 27620 14962 27672 14968
rect 27632 14278 27660 14962
rect 28000 14618 28028 15574
rect 28632 15260 28928 15280
rect 28688 15258 28712 15260
rect 28768 15258 28792 15260
rect 28848 15258 28872 15260
rect 28710 15206 28712 15258
rect 28774 15206 28786 15258
rect 28848 15206 28850 15258
rect 28688 15204 28712 15206
rect 28768 15204 28792 15206
rect 28848 15204 28872 15206
rect 28632 15184 28928 15204
rect 29012 15026 29040 16000
rect 29184 15982 29236 15988
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 30300 14890 30328 17206
rect 30564 17196 30616 17202
rect 30564 17138 30616 17144
rect 30576 16658 30604 17138
rect 30840 17060 30892 17066
rect 30840 17002 30892 17008
rect 30852 16726 30880 17002
rect 30840 16720 30892 16726
rect 30840 16662 30892 16668
rect 30564 16652 30616 16658
rect 30564 16594 30616 16600
rect 30748 16652 30800 16658
rect 30748 16594 30800 16600
rect 30656 16040 30708 16046
rect 30656 15982 30708 15988
rect 29276 14884 29328 14890
rect 29276 14826 29328 14832
rect 30288 14884 30340 14890
rect 30288 14826 30340 14832
rect 29288 14618 29316 14826
rect 27988 14612 28040 14618
rect 27988 14554 28040 14560
rect 29276 14612 29328 14618
rect 29276 14554 29328 14560
rect 27620 14272 27672 14278
rect 27620 14214 27672 14220
rect 26976 13456 27028 13462
rect 26976 13398 27028 13404
rect 26148 13388 26200 13394
rect 26148 13330 26200 13336
rect 26056 12980 26108 12986
rect 26056 12922 26108 12928
rect 26148 12912 26200 12918
rect 26148 12854 26200 12860
rect 25964 12776 26016 12782
rect 25964 12718 26016 12724
rect 25976 12442 26004 12718
rect 25964 12436 26016 12442
rect 25608 12406 25728 12434
rect 25596 12232 25648 12238
rect 25596 12174 25648 12180
rect 25608 11762 25636 12174
rect 25596 11756 25648 11762
rect 25596 11698 25648 11704
rect 25412 11008 25464 11014
rect 25412 10950 25464 10956
rect 25424 10674 25452 10950
rect 25608 10810 25636 11698
rect 25700 11218 25728 12406
rect 25964 12378 26016 12384
rect 25872 12232 25924 12238
rect 25872 12174 25924 12180
rect 25884 11898 25912 12174
rect 25872 11892 25924 11898
rect 25872 11834 25924 11840
rect 25976 11694 26004 12378
rect 26160 12374 26188 12854
rect 27632 12850 27660 14214
rect 28000 13870 28028 14554
rect 28632 14172 28928 14192
rect 28688 14170 28712 14172
rect 28768 14170 28792 14172
rect 28848 14170 28872 14172
rect 28710 14118 28712 14170
rect 28774 14118 28786 14170
rect 28848 14118 28850 14170
rect 28688 14116 28712 14118
rect 28768 14116 28792 14118
rect 28848 14116 28872 14118
rect 28632 14096 28928 14116
rect 27988 13864 28040 13870
rect 27988 13806 28040 13812
rect 28540 13796 28592 13802
rect 28540 13738 28592 13744
rect 28552 13530 28580 13738
rect 29460 13728 29512 13734
rect 29460 13670 29512 13676
rect 28540 13524 28592 13530
rect 28540 13466 28592 13472
rect 28172 13388 28224 13394
rect 28172 13330 28224 13336
rect 28080 13184 28132 13190
rect 28080 13126 28132 13132
rect 28092 12850 28120 13126
rect 26240 12844 26292 12850
rect 26240 12786 26292 12792
rect 27620 12844 27672 12850
rect 27620 12786 27672 12792
rect 27804 12844 27856 12850
rect 27804 12786 27856 12792
rect 28080 12844 28132 12850
rect 28080 12786 28132 12792
rect 26148 12368 26200 12374
rect 26148 12310 26200 12316
rect 26252 11898 26280 12786
rect 27816 12434 27844 12786
rect 27816 12406 27936 12434
rect 26884 12164 26936 12170
rect 26884 12106 26936 12112
rect 26608 12096 26660 12102
rect 26608 12038 26660 12044
rect 26240 11892 26292 11898
rect 26240 11834 26292 11840
rect 26620 11694 26648 12038
rect 25964 11688 26016 11694
rect 25964 11630 26016 11636
rect 26608 11688 26660 11694
rect 26608 11630 26660 11636
rect 26620 11218 26648 11630
rect 26896 11286 26924 12106
rect 27908 11762 27936 12406
rect 27896 11756 27948 11762
rect 27896 11698 27948 11704
rect 27804 11552 27856 11558
rect 27804 11494 27856 11500
rect 27816 11286 27844 11494
rect 26884 11280 26936 11286
rect 26884 11222 26936 11228
rect 27804 11280 27856 11286
rect 27804 11222 27856 11228
rect 25688 11212 25740 11218
rect 25688 11154 25740 11160
rect 26608 11212 26660 11218
rect 26608 11154 26660 11160
rect 25596 10804 25648 10810
rect 25596 10746 25648 10752
rect 25412 10668 25464 10674
rect 25412 10610 25464 10616
rect 25608 10130 25636 10746
rect 25596 10124 25648 10130
rect 25596 10066 25648 10072
rect 25596 5704 25648 5710
rect 25596 5646 25648 5652
rect 25608 5370 25636 5646
rect 25596 5364 25648 5370
rect 25596 5306 25648 5312
rect 25700 5302 25728 11154
rect 25964 11144 26016 11150
rect 25964 11086 26016 11092
rect 25976 9654 26004 11086
rect 26896 10810 26924 11222
rect 27908 11150 27936 11698
rect 28184 11694 28212 13330
rect 28552 12714 28580 13466
rect 28632 13084 28928 13104
rect 28688 13082 28712 13084
rect 28768 13082 28792 13084
rect 28848 13082 28872 13084
rect 28710 13030 28712 13082
rect 28774 13030 28786 13082
rect 28848 13030 28850 13082
rect 28688 13028 28712 13030
rect 28768 13028 28792 13030
rect 28848 13028 28872 13030
rect 28632 13008 28928 13028
rect 28540 12708 28592 12714
rect 28540 12650 28592 12656
rect 28552 12442 28580 12650
rect 28264 12436 28316 12442
rect 28264 12378 28316 12384
rect 28540 12436 28592 12442
rect 28540 12378 28592 12384
rect 28172 11688 28224 11694
rect 28172 11630 28224 11636
rect 27896 11144 27948 11150
rect 27896 11086 27948 11092
rect 26976 11076 27028 11082
rect 26976 11018 27028 11024
rect 26884 10804 26936 10810
rect 26884 10746 26936 10752
rect 25964 9648 26016 9654
rect 25964 9590 26016 9596
rect 25976 9058 26004 9590
rect 25884 9030 26004 9058
rect 25884 7478 25912 9030
rect 25964 8968 26016 8974
rect 25964 8910 26016 8916
rect 25976 8634 26004 8910
rect 26056 8832 26108 8838
rect 26056 8774 26108 8780
rect 25964 8628 26016 8634
rect 25964 8570 26016 8576
rect 26068 8430 26096 8774
rect 26056 8424 26108 8430
rect 26056 8366 26108 8372
rect 25872 7472 25924 7478
rect 25872 7414 25924 7420
rect 26068 7206 26096 8366
rect 26988 7954 27016 11018
rect 27160 10532 27212 10538
rect 27160 10474 27212 10480
rect 27172 10198 27200 10474
rect 27160 10192 27212 10198
rect 27160 10134 27212 10140
rect 27172 10010 27200 10134
rect 27080 9982 27200 10010
rect 27080 9042 27108 9982
rect 27068 9036 27120 9042
rect 27068 8978 27120 8984
rect 26976 7948 27028 7954
rect 26976 7890 27028 7896
rect 27080 7834 27108 8978
rect 28184 8922 28212 11630
rect 28276 11626 28304 12378
rect 29472 12306 29500 13670
rect 30380 13456 30432 13462
rect 30380 13398 30432 13404
rect 29552 13388 29604 13394
rect 29552 13330 29604 13336
rect 29564 12986 29592 13330
rect 29552 12980 29604 12986
rect 29552 12922 29604 12928
rect 30392 12918 30420 13398
rect 30472 13184 30524 13190
rect 30472 13126 30524 13132
rect 30380 12912 30432 12918
rect 30380 12854 30432 12860
rect 29552 12776 29604 12782
rect 29552 12718 29604 12724
rect 29564 12442 29592 12718
rect 30288 12708 30340 12714
rect 30288 12650 30340 12656
rect 29552 12436 29604 12442
rect 30300 12434 30328 12650
rect 29552 12378 29604 12384
rect 30208 12406 30328 12434
rect 29460 12300 29512 12306
rect 29460 12242 29512 12248
rect 28632 11996 28928 12016
rect 28688 11994 28712 11996
rect 28768 11994 28792 11996
rect 28848 11994 28872 11996
rect 28710 11942 28712 11994
rect 28774 11942 28786 11994
rect 28848 11942 28850 11994
rect 28688 11940 28712 11942
rect 28768 11940 28792 11942
rect 28848 11940 28872 11942
rect 28632 11920 28928 11940
rect 28448 11688 28500 11694
rect 28448 11630 28500 11636
rect 29552 11688 29604 11694
rect 29552 11630 29604 11636
rect 28264 11620 28316 11626
rect 28264 11562 28316 11568
rect 28276 11286 28304 11562
rect 28264 11280 28316 11286
rect 28264 11222 28316 11228
rect 28276 10538 28304 11222
rect 28460 11014 28488 11630
rect 29092 11144 29144 11150
rect 29092 11086 29144 11092
rect 28448 11008 28500 11014
rect 28448 10950 28500 10956
rect 28264 10532 28316 10538
rect 28264 10474 28316 10480
rect 28356 9920 28408 9926
rect 28356 9862 28408 9868
rect 28368 9042 28396 9862
rect 28356 9036 28408 9042
rect 28356 8978 28408 8984
rect 28092 8894 28212 8922
rect 27804 7948 27856 7954
rect 27804 7890 27856 7896
rect 26988 7806 27108 7834
rect 26056 7200 26108 7206
rect 26056 7142 26108 7148
rect 26240 7200 26292 7206
rect 26240 7142 26292 7148
rect 25964 6928 26016 6934
rect 26068 6914 26096 7142
rect 26016 6886 26096 6914
rect 25964 6870 26016 6876
rect 26068 6186 26096 6886
rect 26252 6798 26280 7142
rect 26988 6866 27016 7806
rect 27816 6866 27844 7890
rect 28092 7342 28120 8894
rect 28172 8832 28224 8838
rect 28172 8774 28224 8780
rect 28184 8430 28212 8774
rect 28172 8424 28224 8430
rect 28172 8366 28224 8372
rect 28184 7954 28212 8366
rect 28172 7948 28224 7954
rect 28172 7890 28224 7896
rect 28460 7342 28488 10950
rect 28632 10908 28928 10928
rect 28688 10906 28712 10908
rect 28768 10906 28792 10908
rect 28848 10906 28872 10908
rect 28710 10854 28712 10906
rect 28774 10854 28786 10906
rect 28848 10854 28850 10906
rect 28688 10852 28712 10854
rect 28768 10852 28792 10854
rect 28848 10852 28872 10854
rect 28632 10832 28928 10852
rect 29104 10606 29132 11086
rect 29564 10810 29592 11630
rect 29644 11008 29696 11014
rect 29644 10950 29696 10956
rect 29656 10810 29684 10950
rect 29552 10804 29604 10810
rect 29552 10746 29604 10752
rect 29644 10804 29696 10810
rect 29644 10746 29696 10752
rect 29644 10668 29696 10674
rect 29644 10610 29696 10616
rect 29092 10600 29144 10606
rect 29092 10542 29144 10548
rect 29656 10266 29684 10610
rect 29644 10260 29696 10266
rect 29644 10202 29696 10208
rect 29092 9988 29144 9994
rect 29092 9930 29144 9936
rect 28632 9820 28928 9840
rect 28688 9818 28712 9820
rect 28768 9818 28792 9820
rect 28848 9818 28872 9820
rect 28710 9766 28712 9818
rect 28774 9766 28786 9818
rect 28848 9766 28850 9818
rect 28688 9764 28712 9766
rect 28768 9764 28792 9766
rect 28848 9764 28872 9766
rect 28632 9744 28928 9764
rect 29000 9512 29052 9518
rect 29000 9454 29052 9460
rect 28540 8832 28592 8838
rect 28540 8774 28592 8780
rect 28552 8090 28580 8774
rect 28632 8732 28928 8752
rect 28688 8730 28712 8732
rect 28768 8730 28792 8732
rect 28848 8730 28872 8732
rect 28710 8678 28712 8730
rect 28774 8678 28786 8730
rect 28848 8678 28850 8730
rect 28688 8676 28712 8678
rect 28768 8676 28792 8678
rect 28848 8676 28872 8678
rect 28632 8656 28928 8676
rect 28540 8084 28592 8090
rect 28540 8026 28592 8032
rect 28552 7478 28580 8026
rect 29012 8022 29040 9454
rect 29104 9178 29132 9930
rect 29460 9512 29512 9518
rect 29460 9454 29512 9460
rect 29472 9178 29500 9454
rect 29092 9172 29144 9178
rect 29092 9114 29144 9120
rect 29460 9172 29512 9178
rect 29460 9114 29512 9120
rect 29092 8968 29144 8974
rect 29092 8910 29144 8916
rect 29000 8016 29052 8022
rect 29000 7958 29052 7964
rect 28632 7644 28928 7664
rect 28688 7642 28712 7644
rect 28768 7642 28792 7644
rect 28848 7642 28872 7644
rect 28710 7590 28712 7642
rect 28774 7590 28786 7642
rect 28848 7590 28850 7642
rect 28688 7588 28712 7590
rect 28768 7588 28792 7590
rect 28848 7588 28872 7590
rect 28632 7568 28928 7588
rect 28540 7472 28592 7478
rect 28540 7414 28592 7420
rect 29104 7342 29132 8910
rect 29552 8356 29604 8362
rect 29552 8298 29604 8304
rect 29564 8022 29592 8298
rect 29656 8022 29684 10202
rect 30208 10198 30236 12406
rect 30392 12374 30420 12854
rect 30484 12782 30512 13126
rect 30472 12776 30524 12782
rect 30472 12718 30524 12724
rect 30668 12714 30696 15982
rect 30760 15162 30788 16594
rect 30852 15978 30880 16662
rect 30840 15972 30892 15978
rect 30840 15914 30892 15920
rect 30852 15706 30880 15914
rect 30840 15700 30892 15706
rect 30840 15642 30892 15648
rect 30748 15156 30800 15162
rect 30748 15098 30800 15104
rect 30760 14482 30788 15098
rect 30944 14958 30972 18158
rect 31208 17128 31260 17134
rect 31208 17070 31260 17076
rect 31024 16992 31076 16998
rect 31024 16934 31076 16940
rect 31036 16182 31064 16934
rect 31220 16658 31248 17070
rect 31588 16658 31616 18362
rect 31772 17746 31800 19246
rect 32140 18970 32168 19790
rect 32220 19440 32272 19446
rect 32220 19382 32272 19388
rect 32232 19174 32260 19382
rect 32220 19168 32272 19174
rect 32220 19110 32272 19116
rect 32128 18964 32180 18970
rect 32128 18906 32180 18912
rect 32232 18766 32260 19110
rect 32220 18760 32272 18766
rect 32220 18702 32272 18708
rect 31760 17740 31812 17746
rect 31760 17682 31812 17688
rect 32128 17672 32180 17678
rect 32128 17614 32180 17620
rect 32036 17128 32088 17134
rect 32036 17070 32088 17076
rect 31944 16992 31996 16998
rect 31944 16934 31996 16940
rect 31956 16726 31984 16934
rect 31944 16720 31996 16726
rect 31944 16662 31996 16668
rect 31208 16652 31260 16658
rect 31208 16594 31260 16600
rect 31392 16652 31444 16658
rect 31392 16594 31444 16600
rect 31576 16652 31628 16658
rect 31576 16594 31628 16600
rect 31852 16652 31904 16658
rect 31852 16594 31904 16600
rect 31024 16176 31076 16182
rect 31024 16118 31076 16124
rect 31404 16046 31432 16594
rect 31588 16114 31616 16594
rect 31576 16108 31628 16114
rect 31576 16050 31628 16056
rect 31864 16046 31892 16594
rect 32048 16590 32076 17070
rect 32140 16794 32168 17614
rect 32220 17060 32272 17066
rect 32220 17002 32272 17008
rect 32128 16788 32180 16794
rect 32128 16730 32180 16736
rect 32232 16726 32260 17002
rect 32220 16720 32272 16726
rect 32220 16662 32272 16668
rect 32036 16584 32088 16590
rect 32036 16526 32088 16532
rect 31392 16040 31444 16046
rect 31392 15982 31444 15988
rect 31852 16040 31904 16046
rect 31852 15982 31904 15988
rect 31208 15972 31260 15978
rect 31208 15914 31260 15920
rect 31220 15366 31248 15914
rect 31024 15360 31076 15366
rect 31024 15302 31076 15308
rect 31208 15360 31260 15366
rect 31208 15302 31260 15308
rect 30932 14952 30984 14958
rect 30932 14894 30984 14900
rect 30748 14476 30800 14482
rect 30748 14418 30800 14424
rect 30932 13796 30984 13802
rect 30932 13738 30984 13744
rect 30944 12986 30972 13738
rect 31036 13394 31064 15302
rect 31404 14958 31432 15982
rect 32048 15706 32076 16526
rect 32128 15904 32180 15910
rect 32128 15846 32180 15852
rect 32036 15700 32088 15706
rect 32036 15642 32088 15648
rect 31852 15632 31904 15638
rect 31852 15574 31904 15580
rect 31760 15496 31812 15502
rect 31760 15438 31812 15444
rect 31772 15042 31800 15438
rect 31864 15162 31892 15574
rect 31852 15156 31904 15162
rect 31852 15098 31904 15104
rect 31668 15020 31720 15026
rect 31772 15014 31892 15042
rect 31772 15008 31800 15014
rect 31720 14980 31800 15008
rect 31668 14962 31720 14968
rect 31392 14952 31444 14958
rect 31392 14894 31444 14900
rect 31576 14952 31628 14958
rect 31576 14894 31628 14900
rect 31024 13388 31076 13394
rect 31024 13330 31076 13336
rect 30932 12980 30984 12986
rect 30932 12922 30984 12928
rect 30656 12708 30708 12714
rect 30656 12650 30708 12656
rect 31036 12434 31064 13330
rect 31116 12776 31168 12782
rect 31116 12718 31168 12724
rect 30944 12406 31064 12434
rect 30380 12368 30432 12374
rect 30380 12310 30432 12316
rect 30288 12300 30340 12306
rect 30288 12242 30340 12248
rect 30748 12300 30800 12306
rect 30748 12242 30800 12248
rect 30300 12186 30328 12242
rect 30300 12158 30420 12186
rect 30392 11694 30420 12158
rect 30760 11694 30788 12242
rect 30380 11688 30432 11694
rect 30380 11630 30432 11636
rect 30748 11688 30800 11694
rect 30748 11630 30800 11636
rect 30392 10674 30420 11630
rect 30656 11008 30708 11014
rect 30656 10950 30708 10956
rect 30380 10668 30432 10674
rect 30380 10610 30432 10616
rect 30668 10606 30696 10950
rect 30656 10600 30708 10606
rect 30656 10542 30708 10548
rect 30196 10192 30248 10198
rect 30196 10134 30248 10140
rect 29736 9512 29788 9518
rect 29736 9454 29788 9460
rect 29552 8016 29604 8022
rect 29552 7958 29604 7964
rect 29644 8016 29696 8022
rect 29644 7958 29696 7964
rect 29276 7948 29328 7954
rect 29328 7908 29408 7936
rect 29276 7890 29328 7896
rect 28080 7336 28132 7342
rect 28080 7278 28132 7284
rect 28448 7336 28500 7342
rect 28448 7278 28500 7284
rect 29092 7336 29144 7342
rect 29092 7278 29144 7284
rect 26976 6860 27028 6866
rect 26976 6802 27028 6808
rect 27804 6860 27856 6866
rect 27804 6802 27856 6808
rect 26240 6792 26292 6798
rect 26240 6734 26292 6740
rect 26056 6180 26108 6186
rect 26056 6122 26108 6128
rect 25964 6112 26016 6118
rect 25964 6054 26016 6060
rect 25688 5296 25740 5302
rect 25688 5238 25740 5244
rect 25700 4622 25728 5238
rect 25976 5234 26004 6054
rect 26068 5710 26096 6122
rect 26988 5914 27016 6802
rect 28092 6254 28120 7278
rect 28264 6656 28316 6662
rect 28264 6598 28316 6604
rect 28276 6254 28304 6598
rect 28460 6254 28488 7278
rect 28724 7268 28776 7274
rect 28724 7210 28776 7216
rect 28736 7002 28764 7210
rect 28724 6996 28776 7002
rect 28724 6938 28776 6944
rect 28632 6556 28928 6576
rect 28688 6554 28712 6556
rect 28768 6554 28792 6556
rect 28848 6554 28872 6556
rect 28710 6502 28712 6554
rect 28774 6502 28786 6554
rect 28848 6502 28850 6554
rect 28688 6500 28712 6502
rect 28768 6500 28792 6502
rect 28848 6500 28872 6502
rect 28632 6480 28928 6500
rect 28080 6248 28132 6254
rect 28080 6190 28132 6196
rect 28264 6248 28316 6254
rect 28264 6190 28316 6196
rect 28448 6248 28500 6254
rect 28448 6190 28500 6196
rect 27804 6112 27856 6118
rect 27804 6054 27856 6060
rect 26976 5908 27028 5914
rect 26976 5850 27028 5856
rect 27528 5908 27580 5914
rect 27528 5850 27580 5856
rect 26056 5704 26108 5710
rect 26056 5646 26108 5652
rect 26068 5574 26096 5646
rect 26056 5568 26108 5574
rect 26056 5510 26108 5516
rect 27068 5568 27120 5574
rect 27068 5510 27120 5516
rect 25964 5228 26016 5234
rect 25964 5170 26016 5176
rect 27080 5030 27108 5510
rect 27068 5024 27120 5030
rect 27068 4966 27120 4972
rect 25688 4616 25740 4622
rect 25688 4558 25740 4564
rect 27080 4554 27108 4966
rect 27068 4548 27120 4554
rect 27068 4490 27120 4496
rect 26792 4480 26844 4486
rect 26792 4422 26844 4428
rect 26804 3670 26832 4422
rect 27540 4078 27568 5850
rect 27816 5846 27844 6054
rect 27804 5840 27856 5846
rect 27804 5782 27856 5788
rect 28092 4758 28120 6190
rect 28080 4752 28132 4758
rect 28080 4694 28132 4700
rect 28460 4690 28488 6190
rect 29104 5574 29132 7278
rect 29380 6866 29408 7908
rect 29564 7342 29592 7958
rect 29552 7336 29604 7342
rect 29552 7278 29604 7284
rect 29276 6860 29328 6866
rect 29276 6802 29328 6808
rect 29368 6860 29420 6866
rect 29368 6802 29420 6808
rect 29288 6458 29316 6802
rect 29380 6458 29408 6802
rect 29276 6452 29328 6458
rect 29276 6394 29328 6400
rect 29368 6452 29420 6458
rect 29368 6394 29420 6400
rect 29276 6316 29328 6322
rect 29276 6258 29328 6264
rect 29288 5914 29316 6258
rect 29656 6186 29684 7958
rect 29748 7274 29776 9454
rect 30208 8430 30236 10134
rect 30760 10130 30788 11630
rect 30748 10124 30800 10130
rect 30748 10066 30800 10072
rect 30760 9654 30788 10066
rect 30748 9648 30800 9654
rect 30748 9590 30800 9596
rect 30748 9512 30800 9518
rect 30748 9454 30800 9460
rect 30760 9110 30788 9454
rect 30748 9104 30800 9110
rect 30748 9046 30800 9052
rect 30944 9042 30972 12406
rect 31128 12306 31156 12718
rect 31300 12708 31352 12714
rect 31300 12650 31352 12656
rect 31024 12300 31076 12306
rect 31024 12242 31076 12248
rect 31116 12300 31168 12306
rect 31116 12242 31168 12248
rect 31036 11694 31064 12242
rect 31312 11694 31340 12650
rect 31588 12434 31616 14894
rect 31760 14884 31812 14890
rect 31760 14826 31812 14832
rect 31772 13802 31800 14826
rect 31760 13796 31812 13802
rect 31760 13738 31812 13744
rect 31772 12782 31800 13738
rect 31864 13734 31892 15014
rect 32140 14958 32168 15846
rect 32128 14952 32180 14958
rect 32128 14894 32180 14900
rect 32220 14816 32272 14822
rect 32220 14758 32272 14764
rect 32036 14544 32088 14550
rect 32036 14486 32088 14492
rect 31944 14476 31996 14482
rect 31944 14418 31996 14424
rect 31956 13870 31984 14418
rect 31944 13864 31996 13870
rect 31944 13806 31996 13812
rect 31852 13728 31904 13734
rect 31852 13670 31904 13676
rect 31864 13326 31892 13670
rect 31852 13320 31904 13326
rect 31852 13262 31904 13268
rect 31760 12776 31812 12782
rect 31760 12718 31812 12724
rect 31496 12406 31616 12434
rect 31392 11756 31444 11762
rect 31392 11698 31444 11704
rect 31024 11688 31076 11694
rect 31024 11630 31076 11636
rect 31300 11688 31352 11694
rect 31300 11630 31352 11636
rect 31404 11642 31432 11698
rect 31496 11642 31524 12406
rect 31036 11354 31064 11630
rect 31404 11614 31524 11642
rect 31024 11348 31076 11354
rect 31024 11290 31076 11296
rect 31036 10674 31064 11290
rect 31208 11212 31260 11218
rect 31208 11154 31260 11160
rect 31220 10742 31248 11154
rect 31208 10736 31260 10742
rect 31208 10678 31260 10684
rect 31024 10668 31076 10674
rect 31024 10610 31076 10616
rect 31116 10124 31168 10130
rect 31116 10066 31168 10072
rect 30932 9036 30984 9042
rect 30932 8978 30984 8984
rect 30470 8936 30526 8945
rect 30470 8871 30526 8880
rect 30484 8498 30512 8871
rect 30944 8498 30972 8978
rect 31024 8968 31076 8974
rect 31024 8910 31076 8916
rect 30472 8492 30524 8498
rect 30472 8434 30524 8440
rect 30932 8492 30984 8498
rect 30932 8434 30984 8440
rect 29920 8424 29972 8430
rect 29920 8366 29972 8372
rect 30104 8424 30156 8430
rect 30104 8366 30156 8372
rect 30196 8424 30248 8430
rect 30196 8366 30248 8372
rect 29932 8090 29960 8366
rect 29920 8084 29972 8090
rect 29920 8026 29972 8032
rect 29932 7970 29960 8026
rect 29840 7942 29960 7970
rect 30012 7948 30064 7954
rect 29840 7478 29868 7942
rect 30012 7890 30064 7896
rect 29920 7880 29972 7886
rect 29920 7822 29972 7828
rect 29932 7546 29960 7822
rect 29920 7540 29972 7546
rect 29920 7482 29972 7488
rect 30024 7478 30052 7890
rect 30116 7818 30144 8366
rect 30104 7812 30156 7818
rect 30104 7754 30156 7760
rect 29828 7472 29880 7478
rect 29828 7414 29880 7420
rect 30012 7472 30064 7478
rect 30012 7414 30064 7420
rect 29736 7268 29788 7274
rect 29736 7210 29788 7216
rect 29748 6186 29776 7210
rect 30024 6866 30052 7414
rect 30472 7404 30524 7410
rect 30472 7346 30524 7352
rect 30012 6860 30064 6866
rect 30012 6802 30064 6808
rect 30484 6254 30512 7346
rect 30564 7336 30616 7342
rect 30564 7278 30616 7284
rect 30576 6458 30604 7278
rect 31036 6798 31064 8910
rect 31128 8430 31156 10066
rect 31220 9518 31248 10678
rect 31496 10606 31524 11614
rect 31864 11218 31892 13262
rect 31956 12306 31984 13806
rect 31944 12300 31996 12306
rect 31944 12242 31996 12248
rect 31852 11212 31904 11218
rect 31852 11154 31904 11160
rect 31484 10600 31536 10606
rect 31484 10542 31536 10548
rect 31300 10464 31352 10470
rect 31300 10406 31352 10412
rect 31312 10062 31340 10406
rect 31496 10130 31524 10542
rect 31668 10532 31720 10538
rect 31668 10474 31720 10480
rect 31484 10124 31536 10130
rect 31484 10066 31536 10072
rect 31300 10056 31352 10062
rect 31300 9998 31352 10004
rect 31312 9518 31340 9998
rect 31680 9994 31708 10474
rect 31668 9988 31720 9994
rect 31668 9930 31720 9936
rect 31208 9512 31260 9518
rect 31208 9454 31260 9460
rect 31300 9512 31352 9518
rect 31300 9454 31352 9460
rect 31116 8424 31168 8430
rect 31116 8366 31168 8372
rect 31312 7954 31340 9454
rect 31392 8424 31444 8430
rect 31392 8366 31444 8372
rect 31576 8424 31628 8430
rect 31576 8366 31628 8372
rect 31116 7948 31168 7954
rect 31116 7890 31168 7896
rect 31300 7948 31352 7954
rect 31300 7890 31352 7896
rect 31128 7410 31156 7890
rect 31208 7880 31260 7886
rect 31208 7822 31260 7828
rect 31116 7404 31168 7410
rect 31116 7346 31168 7352
rect 31220 7342 31248 7822
rect 31208 7336 31260 7342
rect 31208 7278 31260 7284
rect 31300 7336 31352 7342
rect 31300 7278 31352 7284
rect 31024 6792 31076 6798
rect 31024 6734 31076 6740
rect 30564 6452 30616 6458
rect 30616 6412 30788 6440
rect 30564 6394 30616 6400
rect 30472 6248 30524 6254
rect 30472 6190 30524 6196
rect 29644 6180 29696 6186
rect 29644 6122 29696 6128
rect 29736 6180 29788 6186
rect 29736 6122 29788 6128
rect 29276 5908 29328 5914
rect 29276 5850 29328 5856
rect 30380 5840 30432 5846
rect 30380 5782 30432 5788
rect 29092 5568 29144 5574
rect 29092 5510 29144 5516
rect 28632 5468 28928 5488
rect 28688 5466 28712 5468
rect 28768 5466 28792 5468
rect 28848 5466 28872 5468
rect 28710 5414 28712 5466
rect 28774 5414 28786 5466
rect 28848 5414 28850 5466
rect 28688 5412 28712 5414
rect 28768 5412 28792 5414
rect 28848 5412 28872 5414
rect 28632 5392 28928 5412
rect 28540 4752 28592 4758
rect 28540 4694 28592 4700
rect 27620 4684 27672 4690
rect 27620 4626 27672 4632
rect 28448 4684 28500 4690
rect 28448 4626 28500 4632
rect 27632 4282 27660 4626
rect 28460 4282 28488 4626
rect 27620 4276 27672 4282
rect 27620 4218 27672 4224
rect 28448 4276 28500 4282
rect 28448 4218 28500 4224
rect 28552 4162 28580 4694
rect 28632 4380 28928 4400
rect 28688 4378 28712 4380
rect 28768 4378 28792 4380
rect 28848 4378 28872 4380
rect 28710 4326 28712 4378
rect 28774 4326 28786 4378
rect 28848 4326 28850 4378
rect 28688 4324 28712 4326
rect 28768 4324 28792 4326
rect 28848 4324 28872 4326
rect 28632 4304 28928 4324
rect 29104 4214 29132 5510
rect 30392 5166 30420 5782
rect 30380 5160 30432 5166
rect 30380 5102 30432 5108
rect 30564 5024 30616 5030
rect 30564 4966 30616 4972
rect 30576 4690 30604 4966
rect 30760 4690 30788 6412
rect 31312 6186 31340 7278
rect 31404 7206 31432 8366
rect 31484 8356 31536 8362
rect 31484 8298 31536 8304
rect 31392 7200 31444 7206
rect 31392 7142 31444 7148
rect 31300 6180 31352 6186
rect 31300 6122 31352 6128
rect 31312 5302 31340 6122
rect 31496 5846 31524 8298
rect 31588 7886 31616 8366
rect 31576 7880 31628 7886
rect 31576 7822 31628 7828
rect 31576 6792 31628 6798
rect 31576 6734 31628 6740
rect 31484 5840 31536 5846
rect 31484 5782 31536 5788
rect 31588 5710 31616 6734
rect 31680 6254 31708 9930
rect 31852 8968 31904 8974
rect 31852 8910 31904 8916
rect 31864 8634 31892 8910
rect 31852 8628 31904 8634
rect 31852 8570 31904 8576
rect 32048 6914 32076 14486
rect 32232 14482 32260 14758
rect 32220 14476 32272 14482
rect 32220 14418 32272 14424
rect 32232 13870 32260 14418
rect 32220 13864 32272 13870
rect 32220 13806 32272 13812
rect 32232 13530 32260 13806
rect 32220 13524 32272 13530
rect 32220 13466 32272 13472
rect 32128 13320 32180 13326
rect 32128 13262 32180 13268
rect 32140 12986 32168 13262
rect 32128 12980 32180 12986
rect 32128 12922 32180 12928
rect 32128 12096 32180 12102
rect 32128 12038 32180 12044
rect 32140 11286 32168 12038
rect 32324 11830 32352 34886
rect 32404 29232 32456 29238
rect 32404 29174 32456 29180
rect 32416 28694 32444 29174
rect 32404 28688 32456 28694
rect 32404 28630 32456 28636
rect 32508 12442 32536 34886
rect 33600 33448 33652 33454
rect 33598 33416 33600 33425
rect 33652 33416 33654 33425
rect 33598 33351 33654 33360
rect 33416 33312 33468 33318
rect 33416 33254 33468 33260
rect 33428 32978 33456 33254
rect 33416 32972 33468 32978
rect 33416 32914 33468 32920
rect 33508 32768 33560 32774
rect 33508 32710 33560 32716
rect 33520 32570 33548 32710
rect 33508 32564 33560 32570
rect 33508 32506 33560 32512
rect 33598 29336 33654 29345
rect 33598 29271 33654 29280
rect 33612 29102 33640 29271
rect 33600 29096 33652 29102
rect 33600 29038 33652 29044
rect 33508 28416 33560 28422
rect 33508 28358 33560 28364
rect 33520 27674 33548 28358
rect 33508 27668 33560 27674
rect 33508 27610 33560 27616
rect 33324 27600 33376 27606
rect 33324 27542 33376 27548
rect 32588 27328 32640 27334
rect 32588 27270 32640 27276
rect 32600 26450 32628 27270
rect 33232 26988 33284 26994
rect 33232 26930 33284 26936
rect 32956 26784 33008 26790
rect 32956 26726 33008 26732
rect 32588 26444 32640 26450
rect 32588 26386 32640 26392
rect 32968 24750 32996 26726
rect 33244 26586 33272 26930
rect 33232 26580 33284 26586
rect 33232 26522 33284 26528
rect 33048 26444 33100 26450
rect 33048 26386 33100 26392
rect 33060 25838 33088 26386
rect 33048 25832 33100 25838
rect 33048 25774 33100 25780
rect 33140 25152 33192 25158
rect 33140 25094 33192 25100
rect 32956 24744 33008 24750
rect 32956 24686 33008 24692
rect 32588 24336 32640 24342
rect 32588 24278 32640 24284
rect 32600 23186 32628 24278
rect 32864 24200 32916 24206
rect 32864 24142 32916 24148
rect 32876 23322 32904 24142
rect 32864 23316 32916 23322
rect 32864 23258 32916 23264
rect 32956 23316 33008 23322
rect 32956 23258 33008 23264
rect 32588 23180 32640 23186
rect 32588 23122 32640 23128
rect 32600 22506 32628 23122
rect 32588 22500 32640 22506
rect 32588 22442 32640 22448
rect 32600 21078 32628 22442
rect 32968 21554 32996 23258
rect 33048 22092 33100 22098
rect 33048 22034 33100 22040
rect 32956 21548 33008 21554
rect 32956 21490 33008 21496
rect 32588 21072 32640 21078
rect 32588 21014 32640 21020
rect 32600 20330 32628 21014
rect 32588 20324 32640 20330
rect 32588 20266 32640 20272
rect 32600 19990 32628 20266
rect 32588 19984 32640 19990
rect 32588 19926 32640 19932
rect 32600 18902 32628 19926
rect 33060 19174 33088 22034
rect 33048 19168 33100 19174
rect 33048 19110 33100 19116
rect 32588 18896 32640 18902
rect 32588 18838 32640 18844
rect 32600 17814 32628 18838
rect 32588 17808 32640 17814
rect 32588 17750 32640 17756
rect 32600 17270 32628 17750
rect 32588 17264 32640 17270
rect 32588 17206 32640 17212
rect 32600 15638 32628 17206
rect 33152 17134 33180 25094
rect 33244 24750 33272 26522
rect 33336 25362 33364 27542
rect 33520 26518 33548 27610
rect 33508 26512 33560 26518
rect 33508 26454 33560 26460
rect 33520 25838 33548 26454
rect 33508 25832 33560 25838
rect 33508 25774 33560 25780
rect 33324 25356 33376 25362
rect 33324 25298 33376 25304
rect 33508 25356 33560 25362
rect 33508 25298 33560 25304
rect 33336 24818 33364 25298
rect 33520 25265 33548 25298
rect 33506 25256 33562 25265
rect 33506 25191 33562 25200
rect 33324 24812 33376 24818
rect 33324 24754 33376 24760
rect 33232 24744 33284 24750
rect 33232 24686 33284 24692
rect 33600 24064 33652 24070
rect 33600 24006 33652 24012
rect 33612 23322 33640 24006
rect 33600 23316 33652 23322
rect 33600 23258 33652 23264
rect 33600 21480 33652 21486
rect 33600 21422 33652 21428
rect 33416 21344 33468 21350
rect 33416 21286 33468 21292
rect 33428 21146 33456 21286
rect 33612 21185 33640 21422
rect 33598 21176 33654 21185
rect 33416 21140 33468 21146
rect 33598 21111 33654 21120
rect 33416 21082 33468 21088
rect 33600 19712 33652 19718
rect 33600 19654 33652 19660
rect 33612 19378 33640 19654
rect 33600 19372 33652 19378
rect 33600 19314 33652 19320
rect 33612 18970 33640 19314
rect 33600 18964 33652 18970
rect 33600 18906 33652 18912
rect 33508 17536 33560 17542
rect 33508 17478 33560 17484
rect 33140 17128 33192 17134
rect 33140 17070 33192 17076
rect 33520 16658 33548 17478
rect 33598 17096 33654 17105
rect 33598 17031 33600 17040
rect 33652 17031 33654 17040
rect 33600 17002 33652 17008
rect 33508 16652 33560 16658
rect 33508 16594 33560 16600
rect 33600 16040 33652 16046
rect 33600 15982 33652 15988
rect 33612 15706 33640 15982
rect 33600 15700 33652 15706
rect 33600 15642 33652 15648
rect 32588 15632 32640 15638
rect 32588 15574 32640 15580
rect 33232 14476 33284 14482
rect 33232 14418 33284 14424
rect 33244 13870 33272 14418
rect 33324 14272 33376 14278
rect 33324 14214 33376 14220
rect 33232 13864 33284 13870
rect 33232 13806 33284 13812
rect 32588 13456 32640 13462
rect 32588 13398 32640 13404
rect 32496 12436 32548 12442
rect 32496 12378 32548 12384
rect 32312 11824 32364 11830
rect 32312 11766 32364 11772
rect 32600 11286 32628 13398
rect 33244 13258 33272 13806
rect 33232 13252 33284 13258
rect 33232 13194 33284 13200
rect 33140 12368 33192 12374
rect 33140 12310 33192 12316
rect 32956 12232 33008 12238
rect 32956 12174 33008 12180
rect 32128 11280 32180 11286
rect 32128 11222 32180 11228
rect 32588 11280 32640 11286
rect 32588 11222 32640 11228
rect 32312 10192 32364 10198
rect 32312 10134 32364 10140
rect 32324 8974 32352 10134
rect 32404 10124 32456 10130
rect 32404 10066 32456 10072
rect 32416 9586 32444 10066
rect 32404 9580 32456 9586
rect 32404 9522 32456 9528
rect 32588 9104 32640 9110
rect 32588 9046 32640 9052
rect 32312 8968 32364 8974
rect 32312 8910 32364 8916
rect 32324 7954 32352 8910
rect 32312 7948 32364 7954
rect 32312 7890 32364 7896
rect 32404 7880 32456 7886
rect 32404 7822 32456 7828
rect 32416 7546 32444 7822
rect 32404 7540 32456 7546
rect 32404 7482 32456 7488
rect 32600 6934 32628 9046
rect 32968 8362 32996 12174
rect 33152 10810 33180 12310
rect 33244 11830 33272 13194
rect 33336 12782 33364 14214
rect 33416 13728 33468 13734
rect 33416 13670 33468 13676
rect 33324 12776 33376 12782
rect 33324 12718 33376 12724
rect 33428 12714 33456 13670
rect 33598 13016 33654 13025
rect 33598 12951 33654 12960
rect 33416 12708 33468 12714
rect 33416 12650 33468 12656
rect 33232 11824 33284 11830
rect 33232 11766 33284 11772
rect 33232 11688 33284 11694
rect 33232 11630 33284 11636
rect 33244 11014 33272 11630
rect 33324 11552 33376 11558
rect 33324 11494 33376 11500
rect 33232 11008 33284 11014
rect 33232 10950 33284 10956
rect 33140 10804 33192 10810
rect 33140 10746 33192 10752
rect 33244 10606 33272 10950
rect 33232 10600 33284 10606
rect 33232 10542 33284 10548
rect 33336 10010 33364 11494
rect 33428 10674 33456 12650
rect 33508 12436 33560 12442
rect 33508 12378 33560 12384
rect 33416 10668 33468 10674
rect 33416 10610 33468 10616
rect 33520 10554 33548 12378
rect 33612 12374 33640 12951
rect 33600 12368 33652 12374
rect 33600 12310 33652 12316
rect 33244 9982 33364 10010
rect 33428 10526 33548 10554
rect 33428 9994 33456 10526
rect 33416 9988 33468 9994
rect 33140 9920 33192 9926
rect 33140 9862 33192 9868
rect 33152 8362 33180 9862
rect 33244 9178 33272 9982
rect 33416 9930 33468 9936
rect 33324 9920 33376 9926
rect 33324 9862 33376 9868
rect 33232 9172 33284 9178
rect 33232 9114 33284 9120
rect 33244 8498 33272 9114
rect 33232 8492 33284 8498
rect 33232 8434 33284 8440
rect 32956 8356 33008 8362
rect 32956 8298 33008 8304
rect 33140 8356 33192 8362
rect 33140 8298 33192 8304
rect 31772 6886 32076 6914
rect 32588 6928 32640 6934
rect 31668 6248 31720 6254
rect 31668 6190 31720 6196
rect 31668 6112 31720 6118
rect 31668 6054 31720 6060
rect 31576 5704 31628 5710
rect 31576 5646 31628 5652
rect 31300 5296 31352 5302
rect 31300 5238 31352 5244
rect 31484 5092 31536 5098
rect 31484 5034 31536 5040
rect 30564 4684 30616 4690
rect 30564 4626 30616 4632
rect 30748 4684 30800 4690
rect 30748 4626 30800 4632
rect 31208 4684 31260 4690
rect 31208 4626 31260 4632
rect 29460 4616 29512 4622
rect 29460 4558 29512 4564
rect 29472 4282 29500 4558
rect 29460 4276 29512 4282
rect 29460 4218 29512 4224
rect 29092 4208 29144 4214
rect 28552 4134 28672 4162
rect 29092 4150 29144 4156
rect 28644 4078 28672 4134
rect 27528 4072 27580 4078
rect 27528 4014 27580 4020
rect 28540 4072 28592 4078
rect 28540 4014 28592 4020
rect 28632 4072 28684 4078
rect 28632 4014 28684 4020
rect 29104 4026 29132 4150
rect 29472 4078 29500 4218
rect 30760 4214 30788 4626
rect 31220 4282 31248 4626
rect 31208 4276 31260 4282
rect 31208 4218 31260 4224
rect 30748 4208 30800 4214
rect 30668 4156 30748 4162
rect 30668 4150 30800 4156
rect 30668 4134 30788 4150
rect 31496 4146 31524 5034
rect 31484 4140 31536 4146
rect 29460 4072 29512 4078
rect 27540 3670 27568 4014
rect 28448 4004 28500 4010
rect 28448 3946 28500 3952
rect 26792 3664 26844 3670
rect 26792 3606 26844 3612
rect 27528 3664 27580 3670
rect 27528 3606 27580 3612
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 26528 3194 26556 3470
rect 26516 3188 26568 3194
rect 26516 3130 26568 3136
rect 27540 2854 27568 3606
rect 27528 2848 27580 2854
rect 27528 2790 27580 2796
rect 23097 2748 23393 2768
rect 23153 2746 23177 2748
rect 23233 2746 23257 2748
rect 23313 2746 23337 2748
rect 25148 2746 25820 2774
rect 23175 2694 23177 2746
rect 23239 2694 23251 2746
rect 23313 2694 23315 2746
rect 23153 2692 23177 2694
rect 23233 2692 23257 2694
rect 23313 2692 23337 2694
rect 23097 2672 23393 2692
rect 21916 2644 21968 2650
rect 21916 2586 21968 2592
rect 25792 2582 25820 2746
rect 28460 2582 28488 3946
rect 28552 3670 28580 4014
rect 29104 3998 29224 4026
rect 29460 4014 29512 4020
rect 30288 4072 30340 4078
rect 30288 4014 30340 4020
rect 29092 3936 29144 3942
rect 29092 3878 29144 3884
rect 28540 3664 28592 3670
rect 28540 3606 28592 3612
rect 28632 3292 28928 3312
rect 28688 3290 28712 3292
rect 28768 3290 28792 3292
rect 28848 3290 28872 3292
rect 28710 3238 28712 3290
rect 28774 3238 28786 3290
rect 28848 3238 28850 3290
rect 28688 3236 28712 3238
rect 28768 3236 28792 3238
rect 28848 3236 28872 3238
rect 28632 3216 28928 3236
rect 29104 3058 29132 3878
rect 29196 3602 29224 3998
rect 29552 3936 29604 3942
rect 29552 3878 29604 3884
rect 30196 3936 30248 3942
rect 30196 3878 30248 3884
rect 29564 3738 29592 3878
rect 29552 3732 29604 3738
rect 29552 3674 29604 3680
rect 29184 3596 29236 3602
rect 29184 3538 29236 3544
rect 30208 3398 30236 3878
rect 30300 3534 30328 4014
rect 30380 4004 30432 4010
rect 30380 3946 30432 3952
rect 30288 3528 30340 3534
rect 30288 3470 30340 3476
rect 30196 3392 30248 3398
rect 30196 3334 30248 3340
rect 30300 3194 30328 3470
rect 30288 3188 30340 3194
rect 30288 3130 30340 3136
rect 29092 3052 29144 3058
rect 29092 2994 29144 3000
rect 30392 2582 30420 3946
rect 30668 2990 30696 4134
rect 31484 4082 31536 4088
rect 30748 4072 30800 4078
rect 30748 4014 30800 4020
rect 31208 4072 31260 4078
rect 31208 4014 31260 4020
rect 30760 3602 30788 4014
rect 31220 3670 31248 4014
rect 31496 3738 31524 4082
rect 31484 3732 31536 3738
rect 31484 3674 31536 3680
rect 31208 3664 31260 3670
rect 31208 3606 31260 3612
rect 30748 3596 30800 3602
rect 30748 3538 30800 3544
rect 31220 3194 31248 3606
rect 31588 3602 31616 5646
rect 31680 5166 31708 6054
rect 31668 5160 31720 5166
rect 31668 5102 31720 5108
rect 31576 3596 31628 3602
rect 31576 3538 31628 3544
rect 31208 3188 31260 3194
rect 31208 3130 31260 3136
rect 31588 3126 31616 3538
rect 31576 3120 31628 3126
rect 31576 3062 31628 3068
rect 30656 2984 30708 2990
rect 30656 2926 30708 2932
rect 31772 2582 31800 6886
rect 32640 6886 32904 6914
rect 32588 6870 32640 6876
rect 32876 5846 32904 6886
rect 32968 6254 32996 8298
rect 33152 8090 33180 8298
rect 33140 8084 33192 8090
rect 33140 8026 33192 8032
rect 33244 7834 33272 8434
rect 33336 8430 33364 9862
rect 33428 9722 33456 9930
rect 33416 9716 33468 9722
rect 33416 9658 33468 9664
rect 33324 8424 33376 8430
rect 33324 8366 33376 8372
rect 33416 7948 33468 7954
rect 33416 7890 33468 7896
rect 33600 7948 33652 7954
rect 33600 7890 33652 7896
rect 33244 7806 33364 7834
rect 33232 7744 33284 7750
rect 33232 7686 33284 7692
rect 33140 6792 33192 6798
rect 33140 6734 33192 6740
rect 33152 6458 33180 6734
rect 33140 6452 33192 6458
rect 33140 6394 33192 6400
rect 33244 6254 33272 7686
rect 33336 7274 33364 7806
rect 33428 7478 33456 7890
rect 33416 7472 33468 7478
rect 33416 7414 33468 7420
rect 33324 7268 33376 7274
rect 33324 7210 33376 7216
rect 33612 7002 33640 7890
rect 33600 6996 33652 7002
rect 33600 6938 33652 6944
rect 32956 6248 33008 6254
rect 32956 6190 33008 6196
rect 33232 6248 33284 6254
rect 33232 6190 33284 6196
rect 32864 5840 32916 5846
rect 32864 5782 32916 5788
rect 32128 5704 32180 5710
rect 32128 5646 32180 5652
rect 32140 5370 32168 5646
rect 32312 5568 32364 5574
rect 32312 5510 32364 5516
rect 32128 5364 32180 5370
rect 32128 5306 32180 5312
rect 32324 5234 32352 5510
rect 32312 5228 32364 5234
rect 32312 5170 32364 5176
rect 31944 5160 31996 5166
rect 31944 5102 31996 5108
rect 31852 5024 31904 5030
rect 31852 4966 31904 4972
rect 31864 4826 31892 4966
rect 31852 4820 31904 4826
rect 31852 4762 31904 4768
rect 31956 4706 31984 5102
rect 31864 4690 31984 4706
rect 32324 4690 32352 5170
rect 31852 4684 31984 4690
rect 31904 4678 31984 4684
rect 32312 4684 32364 4690
rect 31852 4626 31904 4632
rect 32312 4626 32364 4632
rect 32496 4548 32548 4554
rect 32496 4490 32548 4496
rect 31852 4480 31904 4486
rect 31852 4422 31904 4428
rect 31864 3670 31892 4422
rect 31852 3664 31904 3670
rect 31852 3606 31904 3612
rect 32508 2582 32536 4490
rect 32876 3670 32904 5782
rect 32968 5166 32996 6190
rect 32956 5160 33008 5166
rect 32956 5102 33008 5108
rect 33048 5160 33100 5166
rect 33048 5102 33100 5108
rect 33060 4622 33088 5102
rect 33416 5024 33468 5030
rect 33416 4966 33468 4972
rect 33428 4758 33456 4966
rect 33598 4856 33654 4865
rect 33598 4791 33654 4800
rect 33612 4758 33640 4791
rect 33416 4752 33468 4758
rect 33416 4694 33468 4700
rect 33600 4752 33652 4758
rect 33600 4694 33652 4700
rect 33048 4616 33100 4622
rect 33048 4558 33100 4564
rect 32864 3664 32916 3670
rect 32864 3606 32916 3612
rect 32876 2922 32904 3606
rect 32864 2916 32916 2922
rect 32864 2858 32916 2864
rect 20720 2576 20772 2582
rect 20720 2518 20772 2524
rect 25780 2576 25832 2582
rect 25780 2518 25832 2524
rect 28448 2576 28500 2582
rect 28448 2518 28500 2524
rect 30380 2576 30432 2582
rect 30380 2518 30432 2524
rect 31760 2576 31812 2582
rect 31760 2518 31812 2524
rect 32496 2576 32548 2582
rect 32496 2518 32548 2524
rect 20536 2508 20588 2514
rect 20536 2450 20588 2456
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 19340 2372 19392 2378
rect 19340 2314 19392 2320
rect 22100 2372 22152 2378
rect 22100 2314 22152 2320
rect 24860 2372 24912 2378
rect 24860 2314 24912 2320
rect 27620 2372 27672 2378
rect 27620 2314 27672 2320
rect 30380 2372 30432 2378
rect 30380 2314 30432 2320
rect 31944 2372 31996 2378
rect 31944 2314 31996 2320
rect 32680 2372 32732 2378
rect 32680 2314 32732 2320
rect 16304 2304 16356 2310
rect 16304 2246 16356 2252
rect 16580 2304 16632 2310
rect 16580 2246 16632 2252
rect 16592 800 16620 2246
rect 17562 2204 17858 2224
rect 17618 2202 17642 2204
rect 17698 2202 17722 2204
rect 17778 2202 17802 2204
rect 17640 2150 17642 2202
rect 17704 2150 17716 2202
rect 17778 2150 17780 2202
rect 17618 2148 17642 2150
rect 17698 2148 17722 2150
rect 17778 2148 17802 2150
rect 17562 2128 17858 2148
rect 19352 800 19380 2314
rect 22112 800 22140 2314
rect 24872 800 24900 2314
rect 27632 800 27660 2314
rect 28632 2204 28928 2224
rect 28688 2202 28712 2204
rect 28768 2202 28792 2204
rect 28848 2202 28872 2204
rect 28710 2150 28712 2202
rect 28774 2150 28786 2202
rect 28848 2150 28850 2202
rect 28688 2148 28712 2150
rect 28768 2148 28792 2150
rect 28848 2148 28872 2150
rect 28632 2128 28928 2148
rect 30392 800 30420 2314
rect 478 0 534 800
rect 2778 0 2834 800
rect 5538 0 5594 800
rect 8298 0 8354 800
rect 11058 0 11114 800
rect 13818 0 13874 800
rect 16578 0 16634 800
rect 19338 0 19394 800
rect 22098 0 22154 800
rect 24858 0 24914 800
rect 27618 0 27674 800
rect 30378 0 30434 800
rect 31956 785 31984 2314
rect 32692 800 32720 2314
rect 31942 776 31998 785
rect 31942 711 31998 720
rect 32678 0 32734 800
<< via2 >>
rect 1398 36760 1454 36816
rect 12026 35386 12082 35388
rect 12106 35386 12162 35388
rect 12186 35386 12242 35388
rect 12266 35386 12322 35388
rect 12026 35334 12052 35386
rect 12052 35334 12082 35386
rect 12106 35334 12116 35386
rect 12116 35334 12162 35386
rect 12186 35334 12232 35386
rect 12232 35334 12242 35386
rect 12266 35334 12296 35386
rect 12296 35334 12322 35386
rect 12026 35332 12082 35334
rect 12106 35332 12162 35334
rect 12186 35332 12242 35334
rect 12266 35332 12322 35334
rect 6491 34842 6547 34844
rect 6571 34842 6627 34844
rect 6651 34842 6707 34844
rect 6731 34842 6787 34844
rect 6491 34790 6517 34842
rect 6517 34790 6547 34842
rect 6571 34790 6581 34842
rect 6581 34790 6627 34842
rect 6651 34790 6697 34842
rect 6697 34790 6707 34842
rect 6731 34790 6761 34842
rect 6761 34790 6787 34842
rect 6491 34788 6547 34790
rect 6571 34788 6627 34790
rect 6651 34788 6707 34790
rect 6731 34788 6787 34790
rect 6491 33754 6547 33756
rect 6571 33754 6627 33756
rect 6651 33754 6707 33756
rect 6731 33754 6787 33756
rect 6491 33702 6517 33754
rect 6517 33702 6547 33754
rect 6571 33702 6581 33754
rect 6581 33702 6627 33754
rect 6651 33702 6697 33754
rect 6697 33702 6707 33754
rect 6731 33702 6761 33754
rect 6761 33702 6787 33754
rect 6491 33700 6547 33702
rect 6571 33700 6627 33702
rect 6651 33700 6707 33702
rect 6731 33700 6787 33702
rect 1398 32680 1454 32736
rect 1766 28600 1822 28656
rect 1398 24520 1454 24576
rect 1398 8200 1454 8256
rect 6491 32666 6547 32668
rect 6571 32666 6627 32668
rect 6651 32666 6707 32668
rect 6731 32666 6787 32668
rect 6491 32614 6517 32666
rect 6517 32614 6547 32666
rect 6571 32614 6581 32666
rect 6581 32614 6627 32666
rect 6651 32614 6697 32666
rect 6697 32614 6707 32666
rect 6731 32614 6761 32666
rect 6761 32614 6787 32666
rect 6491 32612 6547 32614
rect 6571 32612 6627 32614
rect 6651 32612 6707 32614
rect 6731 32612 6787 32614
rect 6491 31578 6547 31580
rect 6571 31578 6627 31580
rect 6651 31578 6707 31580
rect 6731 31578 6787 31580
rect 6491 31526 6517 31578
rect 6517 31526 6547 31578
rect 6571 31526 6581 31578
rect 6581 31526 6627 31578
rect 6651 31526 6697 31578
rect 6697 31526 6707 31578
rect 6731 31526 6761 31578
rect 6761 31526 6787 31578
rect 6491 31524 6547 31526
rect 6571 31524 6627 31526
rect 6651 31524 6707 31526
rect 6731 31524 6787 31526
rect 6491 30490 6547 30492
rect 6571 30490 6627 30492
rect 6651 30490 6707 30492
rect 6731 30490 6787 30492
rect 6491 30438 6517 30490
rect 6517 30438 6547 30490
rect 6571 30438 6581 30490
rect 6581 30438 6627 30490
rect 6651 30438 6697 30490
rect 6697 30438 6707 30490
rect 6731 30438 6761 30490
rect 6761 30438 6787 30490
rect 6491 30436 6547 30438
rect 6571 30436 6627 30438
rect 6651 30436 6707 30438
rect 6731 30436 6787 30438
rect 6491 29402 6547 29404
rect 6571 29402 6627 29404
rect 6651 29402 6707 29404
rect 6731 29402 6787 29404
rect 6491 29350 6517 29402
rect 6517 29350 6547 29402
rect 6571 29350 6581 29402
rect 6581 29350 6627 29402
rect 6651 29350 6697 29402
rect 6697 29350 6707 29402
rect 6731 29350 6761 29402
rect 6761 29350 6787 29402
rect 6491 29348 6547 29350
rect 6571 29348 6627 29350
rect 6651 29348 6707 29350
rect 6731 29348 6787 29350
rect 6491 28314 6547 28316
rect 6571 28314 6627 28316
rect 6651 28314 6707 28316
rect 6731 28314 6787 28316
rect 6491 28262 6517 28314
rect 6517 28262 6547 28314
rect 6571 28262 6581 28314
rect 6581 28262 6627 28314
rect 6651 28262 6697 28314
rect 6697 28262 6707 28314
rect 6731 28262 6761 28314
rect 6761 28262 6787 28314
rect 6491 28260 6547 28262
rect 6571 28260 6627 28262
rect 6651 28260 6707 28262
rect 6731 28260 6787 28262
rect 6491 27226 6547 27228
rect 6571 27226 6627 27228
rect 6651 27226 6707 27228
rect 6731 27226 6787 27228
rect 6491 27174 6517 27226
rect 6517 27174 6547 27226
rect 6571 27174 6581 27226
rect 6581 27174 6627 27226
rect 6651 27174 6697 27226
rect 6697 27174 6707 27226
rect 6731 27174 6761 27226
rect 6761 27174 6787 27226
rect 6491 27172 6547 27174
rect 6571 27172 6627 27174
rect 6651 27172 6707 27174
rect 6731 27172 6787 27174
rect 6491 26138 6547 26140
rect 6571 26138 6627 26140
rect 6651 26138 6707 26140
rect 6731 26138 6787 26140
rect 6491 26086 6517 26138
rect 6517 26086 6547 26138
rect 6571 26086 6581 26138
rect 6581 26086 6627 26138
rect 6651 26086 6697 26138
rect 6697 26086 6707 26138
rect 6731 26086 6761 26138
rect 6761 26086 6787 26138
rect 6491 26084 6547 26086
rect 6571 26084 6627 26086
rect 6651 26084 6707 26086
rect 6731 26084 6787 26086
rect 1766 20460 1822 20496
rect 1766 20440 1768 20460
rect 1768 20440 1820 20460
rect 1820 20440 1822 20460
rect 1766 12316 1768 12336
rect 1768 12316 1820 12336
rect 1820 12316 1822 12336
rect 1766 12280 1822 12316
rect 6491 25050 6547 25052
rect 6571 25050 6627 25052
rect 6651 25050 6707 25052
rect 6731 25050 6787 25052
rect 6491 24998 6517 25050
rect 6517 24998 6547 25050
rect 6571 24998 6581 25050
rect 6581 24998 6627 25050
rect 6651 24998 6697 25050
rect 6697 24998 6707 25050
rect 6731 24998 6761 25050
rect 6761 24998 6787 25050
rect 6491 24996 6547 24998
rect 6571 24996 6627 24998
rect 6651 24996 6707 24998
rect 6731 24996 6787 24998
rect 6491 23962 6547 23964
rect 6571 23962 6627 23964
rect 6651 23962 6707 23964
rect 6731 23962 6787 23964
rect 6491 23910 6517 23962
rect 6517 23910 6547 23962
rect 6571 23910 6581 23962
rect 6581 23910 6627 23962
rect 6651 23910 6697 23962
rect 6697 23910 6707 23962
rect 6731 23910 6761 23962
rect 6761 23910 6787 23962
rect 6491 23908 6547 23910
rect 6571 23908 6627 23910
rect 6651 23908 6707 23910
rect 6731 23908 6787 23910
rect 6491 22874 6547 22876
rect 6571 22874 6627 22876
rect 6651 22874 6707 22876
rect 6731 22874 6787 22876
rect 6491 22822 6517 22874
rect 6517 22822 6547 22874
rect 6571 22822 6581 22874
rect 6581 22822 6627 22874
rect 6651 22822 6697 22874
rect 6697 22822 6707 22874
rect 6731 22822 6761 22874
rect 6761 22822 6787 22874
rect 6491 22820 6547 22822
rect 6571 22820 6627 22822
rect 6651 22820 6707 22822
rect 6731 22820 6787 22822
rect 6491 21786 6547 21788
rect 6571 21786 6627 21788
rect 6651 21786 6707 21788
rect 6731 21786 6787 21788
rect 6491 21734 6517 21786
rect 6517 21734 6547 21786
rect 6571 21734 6581 21786
rect 6581 21734 6627 21786
rect 6651 21734 6697 21786
rect 6697 21734 6707 21786
rect 6731 21734 6761 21786
rect 6761 21734 6787 21786
rect 6491 21732 6547 21734
rect 6571 21732 6627 21734
rect 6651 21732 6707 21734
rect 6731 21732 6787 21734
rect 4066 16360 4122 16416
rect 6491 20698 6547 20700
rect 6571 20698 6627 20700
rect 6651 20698 6707 20700
rect 6731 20698 6787 20700
rect 6491 20646 6517 20698
rect 6517 20646 6547 20698
rect 6571 20646 6581 20698
rect 6581 20646 6627 20698
rect 6651 20646 6697 20698
rect 6697 20646 6707 20698
rect 6731 20646 6761 20698
rect 6761 20646 6787 20698
rect 6491 20644 6547 20646
rect 6571 20644 6627 20646
rect 6651 20644 6707 20646
rect 6731 20644 6787 20646
rect 12026 34298 12082 34300
rect 12106 34298 12162 34300
rect 12186 34298 12242 34300
rect 12266 34298 12322 34300
rect 12026 34246 12052 34298
rect 12052 34246 12082 34298
rect 12106 34246 12116 34298
rect 12116 34246 12162 34298
rect 12186 34246 12232 34298
rect 12232 34246 12242 34298
rect 12266 34246 12296 34298
rect 12296 34246 12322 34298
rect 12026 34244 12082 34246
rect 12106 34244 12162 34246
rect 12186 34244 12242 34246
rect 12266 34244 12322 34246
rect 12026 33210 12082 33212
rect 12106 33210 12162 33212
rect 12186 33210 12242 33212
rect 12266 33210 12322 33212
rect 12026 33158 12052 33210
rect 12052 33158 12082 33210
rect 12106 33158 12116 33210
rect 12116 33158 12162 33210
rect 12186 33158 12232 33210
rect 12232 33158 12242 33210
rect 12266 33158 12296 33210
rect 12296 33158 12322 33210
rect 12026 33156 12082 33158
rect 12106 33156 12162 33158
rect 12186 33156 12242 33158
rect 12266 33156 12322 33158
rect 6491 19610 6547 19612
rect 6571 19610 6627 19612
rect 6651 19610 6707 19612
rect 6731 19610 6787 19612
rect 6491 19558 6517 19610
rect 6517 19558 6547 19610
rect 6571 19558 6581 19610
rect 6581 19558 6627 19610
rect 6651 19558 6697 19610
rect 6697 19558 6707 19610
rect 6731 19558 6761 19610
rect 6761 19558 6787 19610
rect 6491 19556 6547 19558
rect 6571 19556 6627 19558
rect 6651 19556 6707 19558
rect 6731 19556 6787 19558
rect 6491 18522 6547 18524
rect 6571 18522 6627 18524
rect 6651 18522 6707 18524
rect 6731 18522 6787 18524
rect 6491 18470 6517 18522
rect 6517 18470 6547 18522
rect 6571 18470 6581 18522
rect 6581 18470 6627 18522
rect 6651 18470 6697 18522
rect 6697 18470 6707 18522
rect 6731 18470 6761 18522
rect 6761 18470 6787 18522
rect 6491 18468 6547 18470
rect 6571 18468 6627 18470
rect 6651 18468 6707 18470
rect 6731 18468 6787 18470
rect 12026 32122 12082 32124
rect 12106 32122 12162 32124
rect 12186 32122 12242 32124
rect 12266 32122 12322 32124
rect 12026 32070 12052 32122
rect 12052 32070 12082 32122
rect 12106 32070 12116 32122
rect 12116 32070 12162 32122
rect 12186 32070 12232 32122
rect 12232 32070 12242 32122
rect 12266 32070 12296 32122
rect 12296 32070 12322 32122
rect 12026 32068 12082 32070
rect 12106 32068 12162 32070
rect 12186 32068 12242 32070
rect 12266 32068 12322 32070
rect 12026 31034 12082 31036
rect 12106 31034 12162 31036
rect 12186 31034 12242 31036
rect 12266 31034 12322 31036
rect 12026 30982 12052 31034
rect 12052 30982 12082 31034
rect 12106 30982 12116 31034
rect 12116 30982 12162 31034
rect 12186 30982 12232 31034
rect 12232 30982 12242 31034
rect 12266 30982 12296 31034
rect 12296 30982 12322 31034
rect 12026 30980 12082 30982
rect 12106 30980 12162 30982
rect 12186 30980 12242 30982
rect 12266 30980 12322 30982
rect 12026 29946 12082 29948
rect 12106 29946 12162 29948
rect 12186 29946 12242 29948
rect 12266 29946 12322 29948
rect 12026 29894 12052 29946
rect 12052 29894 12082 29946
rect 12106 29894 12116 29946
rect 12116 29894 12162 29946
rect 12186 29894 12232 29946
rect 12232 29894 12242 29946
rect 12266 29894 12296 29946
rect 12296 29894 12322 29946
rect 12026 29892 12082 29894
rect 12106 29892 12162 29894
rect 12186 29892 12242 29894
rect 12266 29892 12322 29894
rect 11150 25356 11206 25392
rect 12026 28858 12082 28860
rect 12106 28858 12162 28860
rect 12186 28858 12242 28860
rect 12266 28858 12322 28860
rect 12026 28806 12052 28858
rect 12052 28806 12082 28858
rect 12106 28806 12116 28858
rect 12116 28806 12162 28858
rect 12186 28806 12232 28858
rect 12232 28806 12242 28858
rect 12266 28806 12296 28858
rect 12296 28806 12322 28858
rect 12026 28804 12082 28806
rect 12106 28804 12162 28806
rect 12186 28804 12242 28806
rect 12266 28804 12322 28806
rect 12026 27770 12082 27772
rect 12106 27770 12162 27772
rect 12186 27770 12242 27772
rect 12266 27770 12322 27772
rect 12026 27718 12052 27770
rect 12052 27718 12082 27770
rect 12106 27718 12116 27770
rect 12116 27718 12162 27770
rect 12186 27718 12232 27770
rect 12232 27718 12242 27770
rect 12266 27718 12296 27770
rect 12296 27718 12322 27770
rect 12026 27716 12082 27718
rect 12106 27716 12162 27718
rect 12186 27716 12242 27718
rect 12266 27716 12322 27718
rect 12026 26682 12082 26684
rect 12106 26682 12162 26684
rect 12186 26682 12242 26684
rect 12266 26682 12322 26684
rect 12026 26630 12052 26682
rect 12052 26630 12082 26682
rect 12106 26630 12116 26682
rect 12116 26630 12162 26682
rect 12186 26630 12232 26682
rect 12232 26630 12242 26682
rect 12266 26630 12296 26682
rect 12296 26630 12322 26682
rect 12026 26628 12082 26630
rect 12106 26628 12162 26630
rect 12186 26628 12242 26630
rect 12266 26628 12322 26630
rect 11150 25336 11152 25356
rect 11152 25336 11204 25356
rect 11204 25336 11206 25356
rect 12026 25594 12082 25596
rect 12106 25594 12162 25596
rect 12186 25594 12242 25596
rect 12266 25594 12322 25596
rect 12026 25542 12052 25594
rect 12052 25542 12082 25594
rect 12106 25542 12116 25594
rect 12116 25542 12162 25594
rect 12186 25542 12232 25594
rect 12232 25542 12242 25594
rect 12266 25542 12296 25594
rect 12296 25542 12322 25594
rect 12026 25540 12082 25542
rect 12106 25540 12162 25542
rect 12186 25540 12242 25542
rect 12266 25540 12322 25542
rect 12026 24506 12082 24508
rect 12106 24506 12162 24508
rect 12186 24506 12242 24508
rect 12266 24506 12322 24508
rect 12026 24454 12052 24506
rect 12052 24454 12082 24506
rect 12106 24454 12116 24506
rect 12116 24454 12162 24506
rect 12186 24454 12232 24506
rect 12232 24454 12242 24506
rect 12266 24454 12296 24506
rect 12296 24454 12322 24506
rect 12026 24452 12082 24454
rect 12106 24452 12162 24454
rect 12186 24452 12242 24454
rect 12266 24452 12322 24454
rect 12026 23418 12082 23420
rect 12106 23418 12162 23420
rect 12186 23418 12242 23420
rect 12266 23418 12322 23420
rect 12026 23366 12052 23418
rect 12052 23366 12082 23418
rect 12106 23366 12116 23418
rect 12116 23366 12162 23418
rect 12186 23366 12232 23418
rect 12232 23366 12242 23418
rect 12266 23366 12296 23418
rect 12296 23366 12322 23418
rect 12026 23364 12082 23366
rect 12106 23364 12162 23366
rect 12186 23364 12242 23366
rect 12266 23364 12322 23366
rect 6491 17434 6547 17436
rect 6571 17434 6627 17436
rect 6651 17434 6707 17436
rect 6731 17434 6787 17436
rect 6491 17382 6517 17434
rect 6517 17382 6547 17434
rect 6571 17382 6581 17434
rect 6581 17382 6627 17434
rect 6651 17382 6697 17434
rect 6697 17382 6707 17434
rect 6731 17382 6761 17434
rect 6761 17382 6787 17434
rect 6491 17380 6547 17382
rect 6571 17380 6627 17382
rect 6651 17380 6707 17382
rect 6731 17380 6787 17382
rect 6491 16346 6547 16348
rect 6571 16346 6627 16348
rect 6651 16346 6707 16348
rect 6731 16346 6787 16348
rect 6491 16294 6517 16346
rect 6517 16294 6547 16346
rect 6571 16294 6581 16346
rect 6581 16294 6627 16346
rect 6651 16294 6697 16346
rect 6697 16294 6707 16346
rect 6731 16294 6761 16346
rect 6761 16294 6787 16346
rect 6491 16292 6547 16294
rect 6571 16292 6627 16294
rect 6651 16292 6707 16294
rect 6731 16292 6787 16294
rect 6491 15258 6547 15260
rect 6571 15258 6627 15260
rect 6651 15258 6707 15260
rect 6731 15258 6787 15260
rect 6491 15206 6517 15258
rect 6517 15206 6547 15258
rect 6571 15206 6581 15258
rect 6581 15206 6627 15258
rect 6651 15206 6697 15258
rect 6697 15206 6707 15258
rect 6731 15206 6761 15258
rect 6761 15206 6787 15258
rect 6491 15204 6547 15206
rect 6571 15204 6627 15206
rect 6651 15204 6707 15206
rect 6731 15204 6787 15206
rect 6491 14170 6547 14172
rect 6571 14170 6627 14172
rect 6651 14170 6707 14172
rect 6731 14170 6787 14172
rect 6491 14118 6517 14170
rect 6517 14118 6547 14170
rect 6571 14118 6581 14170
rect 6581 14118 6627 14170
rect 6651 14118 6697 14170
rect 6697 14118 6707 14170
rect 6731 14118 6761 14170
rect 6761 14118 6787 14170
rect 6491 14116 6547 14118
rect 6571 14116 6627 14118
rect 6651 14116 6707 14118
rect 6731 14116 6787 14118
rect 6491 13082 6547 13084
rect 6571 13082 6627 13084
rect 6651 13082 6707 13084
rect 6731 13082 6787 13084
rect 6491 13030 6517 13082
rect 6517 13030 6547 13082
rect 6571 13030 6581 13082
rect 6581 13030 6627 13082
rect 6651 13030 6697 13082
rect 6697 13030 6707 13082
rect 6731 13030 6761 13082
rect 6761 13030 6787 13082
rect 6491 13028 6547 13030
rect 6571 13028 6627 13030
rect 6651 13028 6707 13030
rect 6731 13028 6787 13030
rect 6491 11994 6547 11996
rect 6571 11994 6627 11996
rect 6651 11994 6707 11996
rect 6731 11994 6787 11996
rect 6491 11942 6517 11994
rect 6517 11942 6547 11994
rect 6571 11942 6581 11994
rect 6581 11942 6627 11994
rect 6651 11942 6697 11994
rect 6697 11942 6707 11994
rect 6731 11942 6761 11994
rect 6761 11942 6787 11994
rect 6491 11940 6547 11942
rect 6571 11940 6627 11942
rect 6651 11940 6707 11942
rect 6731 11940 6787 11942
rect 12026 22330 12082 22332
rect 12106 22330 12162 22332
rect 12186 22330 12242 22332
rect 12266 22330 12322 22332
rect 12026 22278 12052 22330
rect 12052 22278 12082 22330
rect 12106 22278 12116 22330
rect 12116 22278 12162 22330
rect 12186 22278 12232 22330
rect 12232 22278 12242 22330
rect 12266 22278 12296 22330
rect 12296 22278 12322 22330
rect 12026 22276 12082 22278
rect 12106 22276 12162 22278
rect 12186 22276 12242 22278
rect 12266 22276 12322 22278
rect 12162 21956 12218 21992
rect 12162 21936 12164 21956
rect 12164 21936 12216 21956
rect 12216 21936 12218 21956
rect 12026 21242 12082 21244
rect 12106 21242 12162 21244
rect 12186 21242 12242 21244
rect 12266 21242 12322 21244
rect 12026 21190 12052 21242
rect 12052 21190 12082 21242
rect 12106 21190 12116 21242
rect 12116 21190 12162 21242
rect 12186 21190 12232 21242
rect 12232 21190 12242 21242
rect 12266 21190 12296 21242
rect 12296 21190 12322 21242
rect 12026 21188 12082 21190
rect 12106 21188 12162 21190
rect 12186 21188 12242 21190
rect 12266 21188 12322 21190
rect 12806 25372 12808 25392
rect 12808 25372 12860 25392
rect 12860 25372 12862 25392
rect 12806 25336 12862 25372
rect 12026 20154 12082 20156
rect 12106 20154 12162 20156
rect 12186 20154 12242 20156
rect 12266 20154 12322 20156
rect 12026 20102 12052 20154
rect 12052 20102 12082 20154
rect 12106 20102 12116 20154
rect 12116 20102 12162 20154
rect 12186 20102 12232 20154
rect 12232 20102 12242 20154
rect 12266 20102 12296 20154
rect 12296 20102 12322 20154
rect 12026 20100 12082 20102
rect 12106 20100 12162 20102
rect 12186 20100 12242 20102
rect 12266 20100 12322 20102
rect 6491 10906 6547 10908
rect 6571 10906 6627 10908
rect 6651 10906 6707 10908
rect 6731 10906 6787 10908
rect 6491 10854 6517 10906
rect 6517 10854 6547 10906
rect 6571 10854 6581 10906
rect 6581 10854 6627 10906
rect 6651 10854 6697 10906
rect 6697 10854 6707 10906
rect 6731 10854 6761 10906
rect 6761 10854 6787 10906
rect 6491 10852 6547 10854
rect 6571 10852 6627 10854
rect 6651 10852 6707 10854
rect 6731 10852 6787 10854
rect 6491 9818 6547 9820
rect 6571 9818 6627 9820
rect 6651 9818 6707 9820
rect 6731 9818 6787 9820
rect 6491 9766 6517 9818
rect 6517 9766 6547 9818
rect 6571 9766 6581 9818
rect 6581 9766 6627 9818
rect 6651 9766 6697 9818
rect 6697 9766 6707 9818
rect 6731 9766 6761 9818
rect 6761 9766 6787 9818
rect 6491 9764 6547 9766
rect 6571 9764 6627 9766
rect 6651 9764 6707 9766
rect 6731 9764 6787 9766
rect 6491 8730 6547 8732
rect 6571 8730 6627 8732
rect 6651 8730 6707 8732
rect 6731 8730 6787 8732
rect 6491 8678 6517 8730
rect 6517 8678 6547 8730
rect 6571 8678 6581 8730
rect 6581 8678 6627 8730
rect 6651 8678 6697 8730
rect 6697 8678 6707 8730
rect 6731 8678 6761 8730
rect 6761 8678 6787 8730
rect 6491 8676 6547 8678
rect 6571 8676 6627 8678
rect 6651 8676 6707 8678
rect 6731 8676 6787 8678
rect 1858 4120 1914 4176
rect 6491 7642 6547 7644
rect 6571 7642 6627 7644
rect 6651 7642 6707 7644
rect 6731 7642 6787 7644
rect 6491 7590 6517 7642
rect 6517 7590 6547 7642
rect 6571 7590 6581 7642
rect 6581 7590 6627 7642
rect 6651 7590 6697 7642
rect 6697 7590 6707 7642
rect 6731 7590 6761 7642
rect 6761 7590 6787 7642
rect 6491 7588 6547 7590
rect 6571 7588 6627 7590
rect 6651 7588 6707 7590
rect 6731 7588 6787 7590
rect 6491 6554 6547 6556
rect 6571 6554 6627 6556
rect 6651 6554 6707 6556
rect 6731 6554 6787 6556
rect 6491 6502 6517 6554
rect 6517 6502 6547 6554
rect 6571 6502 6581 6554
rect 6581 6502 6627 6554
rect 6651 6502 6697 6554
rect 6697 6502 6707 6554
rect 6731 6502 6761 6554
rect 6761 6502 6787 6554
rect 6491 6500 6547 6502
rect 6571 6500 6627 6502
rect 6651 6500 6707 6502
rect 6731 6500 6787 6502
rect 6491 5466 6547 5468
rect 6571 5466 6627 5468
rect 6651 5466 6707 5468
rect 6731 5466 6787 5468
rect 6491 5414 6517 5466
rect 6517 5414 6547 5466
rect 6571 5414 6581 5466
rect 6581 5414 6627 5466
rect 6651 5414 6697 5466
rect 6697 5414 6707 5466
rect 6731 5414 6761 5466
rect 6761 5414 6787 5466
rect 6491 5412 6547 5414
rect 6571 5412 6627 5414
rect 6651 5412 6707 5414
rect 6731 5412 6787 5414
rect 6491 4378 6547 4380
rect 6571 4378 6627 4380
rect 6651 4378 6707 4380
rect 6731 4378 6787 4380
rect 6491 4326 6517 4378
rect 6517 4326 6547 4378
rect 6571 4326 6581 4378
rect 6581 4326 6627 4378
rect 6651 4326 6697 4378
rect 6697 4326 6707 4378
rect 6731 4326 6761 4378
rect 6761 4326 6787 4378
rect 6491 4324 6547 4326
rect 6571 4324 6627 4326
rect 6651 4324 6707 4326
rect 6731 4324 6787 4326
rect 6491 3290 6547 3292
rect 6571 3290 6627 3292
rect 6651 3290 6707 3292
rect 6731 3290 6787 3292
rect 6491 3238 6517 3290
rect 6517 3238 6547 3290
rect 6571 3238 6581 3290
rect 6581 3238 6627 3290
rect 6651 3238 6697 3290
rect 6697 3238 6707 3290
rect 6731 3238 6761 3290
rect 6761 3238 6787 3290
rect 6491 3236 6547 3238
rect 6571 3236 6627 3238
rect 6651 3236 6707 3238
rect 6731 3236 6787 3238
rect 12026 19066 12082 19068
rect 12106 19066 12162 19068
rect 12186 19066 12242 19068
rect 12266 19066 12322 19068
rect 12026 19014 12052 19066
rect 12052 19014 12082 19066
rect 12106 19014 12116 19066
rect 12116 19014 12162 19066
rect 12186 19014 12232 19066
rect 12232 19014 12242 19066
rect 12266 19014 12296 19066
rect 12296 19014 12322 19066
rect 12026 19012 12082 19014
rect 12106 19012 12162 19014
rect 12186 19012 12242 19014
rect 12266 19012 12322 19014
rect 12254 18536 12310 18592
rect 12026 17978 12082 17980
rect 12106 17978 12162 17980
rect 12186 17978 12242 17980
rect 12266 17978 12322 17980
rect 12026 17926 12052 17978
rect 12052 17926 12082 17978
rect 12106 17926 12116 17978
rect 12116 17926 12162 17978
rect 12186 17926 12232 17978
rect 12232 17926 12242 17978
rect 12266 17926 12296 17978
rect 12296 17926 12322 17978
rect 12026 17924 12082 17926
rect 12106 17924 12162 17926
rect 12186 17924 12242 17926
rect 12266 17924 12322 17926
rect 12026 16890 12082 16892
rect 12106 16890 12162 16892
rect 12186 16890 12242 16892
rect 12266 16890 12322 16892
rect 12026 16838 12052 16890
rect 12052 16838 12082 16890
rect 12106 16838 12116 16890
rect 12116 16838 12162 16890
rect 12186 16838 12232 16890
rect 12232 16838 12242 16890
rect 12266 16838 12296 16890
rect 12296 16838 12322 16890
rect 12026 16836 12082 16838
rect 12106 16836 12162 16838
rect 12186 16836 12242 16838
rect 12266 16836 12322 16838
rect 12026 15802 12082 15804
rect 12106 15802 12162 15804
rect 12186 15802 12242 15804
rect 12266 15802 12322 15804
rect 12026 15750 12052 15802
rect 12052 15750 12082 15802
rect 12106 15750 12116 15802
rect 12116 15750 12162 15802
rect 12186 15750 12232 15802
rect 12232 15750 12242 15802
rect 12266 15750 12296 15802
rect 12296 15750 12322 15802
rect 12026 15748 12082 15750
rect 12106 15748 12162 15750
rect 12186 15748 12242 15750
rect 12266 15748 12322 15750
rect 13358 19252 13360 19272
rect 13360 19252 13412 19272
rect 13412 19252 13414 19272
rect 13358 19216 13414 19252
rect 12026 14714 12082 14716
rect 12106 14714 12162 14716
rect 12186 14714 12242 14716
rect 12266 14714 12322 14716
rect 12026 14662 12052 14714
rect 12052 14662 12082 14714
rect 12106 14662 12116 14714
rect 12116 14662 12162 14714
rect 12186 14662 12232 14714
rect 12232 14662 12242 14714
rect 12266 14662 12296 14714
rect 12296 14662 12322 14714
rect 12026 14660 12082 14662
rect 12106 14660 12162 14662
rect 12186 14660 12242 14662
rect 12266 14660 12322 14662
rect 12026 13626 12082 13628
rect 12106 13626 12162 13628
rect 12186 13626 12242 13628
rect 12266 13626 12322 13628
rect 12026 13574 12052 13626
rect 12052 13574 12082 13626
rect 12106 13574 12116 13626
rect 12116 13574 12162 13626
rect 12186 13574 12232 13626
rect 12232 13574 12242 13626
rect 12266 13574 12296 13626
rect 12296 13574 12322 13626
rect 12026 13572 12082 13574
rect 12106 13572 12162 13574
rect 12186 13572 12242 13574
rect 12266 13572 12322 13574
rect 12026 12538 12082 12540
rect 12106 12538 12162 12540
rect 12186 12538 12242 12540
rect 12266 12538 12322 12540
rect 12026 12486 12052 12538
rect 12052 12486 12082 12538
rect 12106 12486 12116 12538
rect 12116 12486 12162 12538
rect 12186 12486 12232 12538
rect 12232 12486 12242 12538
rect 12266 12486 12296 12538
rect 12296 12486 12322 12538
rect 12026 12484 12082 12486
rect 12106 12484 12162 12486
rect 12186 12484 12242 12486
rect 12266 12484 12322 12486
rect 12026 11450 12082 11452
rect 12106 11450 12162 11452
rect 12186 11450 12242 11452
rect 12266 11450 12322 11452
rect 12026 11398 12052 11450
rect 12052 11398 12082 11450
rect 12106 11398 12116 11450
rect 12116 11398 12162 11450
rect 12186 11398 12232 11450
rect 12232 11398 12242 11450
rect 12266 11398 12296 11450
rect 12296 11398 12322 11450
rect 12026 11396 12082 11398
rect 12106 11396 12162 11398
rect 12186 11396 12242 11398
rect 12266 11396 12322 11398
rect 12026 10362 12082 10364
rect 12106 10362 12162 10364
rect 12186 10362 12242 10364
rect 12266 10362 12322 10364
rect 12026 10310 12052 10362
rect 12052 10310 12082 10362
rect 12106 10310 12116 10362
rect 12116 10310 12162 10362
rect 12186 10310 12232 10362
rect 12232 10310 12242 10362
rect 12266 10310 12296 10362
rect 12296 10310 12322 10362
rect 12026 10308 12082 10310
rect 12106 10308 12162 10310
rect 12186 10308 12242 10310
rect 12266 10308 12322 10310
rect 12026 9274 12082 9276
rect 12106 9274 12162 9276
rect 12186 9274 12242 9276
rect 12266 9274 12322 9276
rect 12026 9222 12052 9274
rect 12052 9222 12082 9274
rect 12106 9222 12116 9274
rect 12116 9222 12162 9274
rect 12186 9222 12232 9274
rect 12232 9222 12242 9274
rect 12266 9222 12296 9274
rect 12296 9222 12322 9274
rect 12026 9220 12082 9222
rect 12106 9220 12162 9222
rect 12186 9220 12242 9222
rect 12266 9220 12322 9222
rect 12026 8186 12082 8188
rect 12106 8186 12162 8188
rect 12186 8186 12242 8188
rect 12266 8186 12322 8188
rect 12026 8134 12052 8186
rect 12052 8134 12082 8186
rect 12106 8134 12116 8186
rect 12116 8134 12162 8186
rect 12186 8134 12232 8186
rect 12232 8134 12242 8186
rect 12266 8134 12296 8186
rect 12296 8134 12322 8186
rect 12026 8132 12082 8134
rect 12106 8132 12162 8134
rect 12186 8132 12242 8134
rect 12266 8132 12322 8134
rect 12026 7098 12082 7100
rect 12106 7098 12162 7100
rect 12186 7098 12242 7100
rect 12266 7098 12322 7100
rect 12026 7046 12052 7098
rect 12052 7046 12082 7098
rect 12106 7046 12116 7098
rect 12116 7046 12162 7098
rect 12186 7046 12232 7098
rect 12232 7046 12242 7098
rect 12266 7046 12296 7098
rect 12296 7046 12322 7098
rect 12026 7044 12082 7046
rect 12106 7044 12162 7046
rect 12186 7044 12242 7046
rect 12266 7044 12322 7046
rect 12026 6010 12082 6012
rect 12106 6010 12162 6012
rect 12186 6010 12242 6012
rect 12266 6010 12322 6012
rect 12026 5958 12052 6010
rect 12052 5958 12082 6010
rect 12106 5958 12116 6010
rect 12116 5958 12162 6010
rect 12186 5958 12232 6010
rect 12232 5958 12242 6010
rect 12266 5958 12296 6010
rect 12296 5958 12322 6010
rect 12026 5956 12082 5958
rect 12106 5956 12162 5958
rect 12186 5956 12242 5958
rect 12266 5956 12322 5958
rect 12026 4922 12082 4924
rect 12106 4922 12162 4924
rect 12186 4922 12242 4924
rect 12266 4922 12322 4924
rect 12026 4870 12052 4922
rect 12052 4870 12082 4922
rect 12106 4870 12116 4922
rect 12116 4870 12162 4922
rect 12186 4870 12232 4922
rect 12232 4870 12242 4922
rect 12266 4870 12296 4922
rect 12296 4870 12322 4922
rect 12026 4868 12082 4870
rect 12106 4868 12162 4870
rect 12186 4868 12242 4870
rect 12266 4868 12322 4870
rect 12026 3834 12082 3836
rect 12106 3834 12162 3836
rect 12186 3834 12242 3836
rect 12266 3834 12322 3836
rect 12026 3782 12052 3834
rect 12052 3782 12082 3834
rect 12106 3782 12116 3834
rect 12116 3782 12162 3834
rect 12186 3782 12232 3834
rect 12232 3782 12242 3834
rect 12266 3782 12296 3834
rect 12296 3782 12322 3834
rect 12026 3780 12082 3782
rect 12106 3780 12162 3782
rect 12186 3780 12242 3782
rect 12266 3780 12322 3782
rect 12026 2746 12082 2748
rect 12106 2746 12162 2748
rect 12186 2746 12242 2748
rect 12266 2746 12322 2748
rect 12026 2694 12052 2746
rect 12052 2694 12082 2746
rect 12106 2694 12116 2746
rect 12116 2694 12162 2746
rect 12186 2694 12232 2746
rect 12232 2694 12242 2746
rect 12266 2694 12296 2746
rect 12296 2694 12322 2746
rect 12026 2692 12082 2694
rect 12106 2692 12162 2694
rect 12186 2692 12242 2694
rect 12266 2692 12322 2694
rect 14646 19216 14702 19272
rect 23097 35386 23153 35388
rect 23177 35386 23233 35388
rect 23257 35386 23313 35388
rect 23337 35386 23393 35388
rect 23097 35334 23123 35386
rect 23123 35334 23153 35386
rect 23177 35334 23187 35386
rect 23187 35334 23233 35386
rect 23257 35334 23303 35386
rect 23303 35334 23313 35386
rect 23337 35334 23367 35386
rect 23367 35334 23393 35386
rect 23097 35332 23153 35334
rect 23177 35332 23233 35334
rect 23257 35332 23313 35334
rect 23337 35332 23393 35334
rect 17562 34842 17618 34844
rect 17642 34842 17698 34844
rect 17722 34842 17778 34844
rect 17802 34842 17858 34844
rect 17562 34790 17588 34842
rect 17588 34790 17618 34842
rect 17642 34790 17652 34842
rect 17652 34790 17698 34842
rect 17722 34790 17768 34842
rect 17768 34790 17778 34842
rect 17802 34790 17832 34842
rect 17832 34790 17858 34842
rect 17562 34788 17618 34790
rect 17642 34788 17698 34790
rect 17722 34788 17778 34790
rect 17802 34788 17858 34790
rect 17562 33754 17618 33756
rect 17642 33754 17698 33756
rect 17722 33754 17778 33756
rect 17802 33754 17858 33756
rect 17562 33702 17588 33754
rect 17588 33702 17618 33754
rect 17642 33702 17652 33754
rect 17652 33702 17698 33754
rect 17722 33702 17768 33754
rect 17768 33702 17778 33754
rect 17802 33702 17832 33754
rect 17832 33702 17858 33754
rect 17562 33700 17618 33702
rect 17642 33700 17698 33702
rect 17722 33700 17778 33702
rect 17802 33700 17858 33702
rect 17562 32666 17618 32668
rect 17642 32666 17698 32668
rect 17722 32666 17778 32668
rect 17802 32666 17858 32668
rect 17562 32614 17588 32666
rect 17588 32614 17618 32666
rect 17642 32614 17652 32666
rect 17652 32614 17698 32666
rect 17722 32614 17768 32666
rect 17768 32614 17778 32666
rect 17802 32614 17832 32666
rect 17832 32614 17858 32666
rect 17562 32612 17618 32614
rect 17642 32612 17698 32614
rect 17722 32612 17778 32614
rect 17802 32612 17858 32614
rect 17562 31578 17618 31580
rect 17642 31578 17698 31580
rect 17722 31578 17778 31580
rect 17802 31578 17858 31580
rect 17562 31526 17588 31578
rect 17588 31526 17618 31578
rect 17642 31526 17652 31578
rect 17652 31526 17698 31578
rect 17722 31526 17768 31578
rect 17768 31526 17778 31578
rect 17802 31526 17832 31578
rect 17832 31526 17858 31578
rect 17562 31524 17618 31526
rect 17642 31524 17698 31526
rect 17722 31524 17778 31526
rect 17802 31524 17858 31526
rect 17562 30490 17618 30492
rect 17642 30490 17698 30492
rect 17722 30490 17778 30492
rect 17802 30490 17858 30492
rect 17562 30438 17588 30490
rect 17588 30438 17618 30490
rect 17642 30438 17652 30490
rect 17652 30438 17698 30490
rect 17722 30438 17768 30490
rect 17768 30438 17778 30490
rect 17802 30438 17832 30490
rect 17832 30438 17858 30490
rect 17562 30436 17618 30438
rect 17642 30436 17698 30438
rect 17722 30436 17778 30438
rect 17802 30436 17858 30438
rect 17562 29402 17618 29404
rect 17642 29402 17698 29404
rect 17722 29402 17778 29404
rect 17802 29402 17858 29404
rect 17562 29350 17588 29402
rect 17588 29350 17618 29402
rect 17642 29350 17652 29402
rect 17652 29350 17698 29402
rect 17722 29350 17768 29402
rect 17768 29350 17778 29402
rect 17802 29350 17832 29402
rect 17832 29350 17858 29402
rect 17562 29348 17618 29350
rect 17642 29348 17698 29350
rect 17722 29348 17778 29350
rect 17802 29348 17858 29350
rect 17562 28314 17618 28316
rect 17642 28314 17698 28316
rect 17722 28314 17778 28316
rect 17802 28314 17858 28316
rect 17562 28262 17588 28314
rect 17588 28262 17618 28314
rect 17642 28262 17652 28314
rect 17652 28262 17698 28314
rect 17722 28262 17768 28314
rect 17768 28262 17778 28314
rect 17802 28262 17832 28314
rect 17832 28262 17858 28314
rect 17562 28260 17618 28262
rect 17642 28260 17698 28262
rect 17722 28260 17778 28262
rect 17802 28260 17858 28262
rect 17562 27226 17618 27228
rect 17642 27226 17698 27228
rect 17722 27226 17778 27228
rect 17802 27226 17858 27228
rect 17562 27174 17588 27226
rect 17588 27174 17618 27226
rect 17642 27174 17652 27226
rect 17652 27174 17698 27226
rect 17722 27174 17768 27226
rect 17768 27174 17778 27226
rect 17802 27174 17832 27226
rect 17832 27174 17858 27226
rect 17562 27172 17618 27174
rect 17642 27172 17698 27174
rect 17722 27172 17778 27174
rect 17802 27172 17858 27174
rect 17562 26138 17618 26140
rect 17642 26138 17698 26140
rect 17722 26138 17778 26140
rect 17802 26138 17858 26140
rect 17562 26086 17588 26138
rect 17588 26086 17618 26138
rect 17642 26086 17652 26138
rect 17652 26086 17698 26138
rect 17722 26086 17768 26138
rect 17768 26086 17778 26138
rect 17802 26086 17832 26138
rect 17832 26086 17858 26138
rect 17562 26084 17618 26086
rect 17642 26084 17698 26086
rect 17722 26084 17778 26086
rect 17802 26084 17858 26086
rect 17562 25050 17618 25052
rect 17642 25050 17698 25052
rect 17722 25050 17778 25052
rect 17802 25050 17858 25052
rect 17562 24998 17588 25050
rect 17588 24998 17618 25050
rect 17642 24998 17652 25050
rect 17652 24998 17698 25050
rect 17722 24998 17768 25050
rect 17768 24998 17778 25050
rect 17802 24998 17832 25050
rect 17832 24998 17858 25050
rect 17562 24996 17618 24998
rect 17642 24996 17698 24998
rect 17722 24996 17778 24998
rect 17802 24996 17858 24998
rect 17562 23962 17618 23964
rect 17642 23962 17698 23964
rect 17722 23962 17778 23964
rect 17802 23962 17858 23964
rect 17562 23910 17588 23962
rect 17588 23910 17618 23962
rect 17642 23910 17652 23962
rect 17652 23910 17698 23962
rect 17722 23910 17768 23962
rect 17768 23910 17778 23962
rect 17802 23910 17832 23962
rect 17832 23910 17858 23962
rect 17562 23908 17618 23910
rect 17642 23908 17698 23910
rect 17722 23908 17778 23910
rect 17802 23908 17858 23910
rect 15014 19236 15070 19272
rect 15014 19216 15016 19236
rect 15016 19216 15068 19236
rect 15068 19216 15070 19236
rect 16578 21936 16634 21992
rect 17562 22874 17618 22876
rect 17642 22874 17698 22876
rect 17722 22874 17778 22876
rect 17802 22874 17858 22876
rect 17562 22822 17588 22874
rect 17588 22822 17618 22874
rect 17642 22822 17652 22874
rect 17652 22822 17698 22874
rect 17722 22822 17768 22874
rect 17768 22822 17778 22874
rect 17802 22822 17832 22874
rect 17832 22822 17858 22874
rect 17562 22820 17618 22822
rect 17642 22820 17698 22822
rect 17722 22820 17778 22822
rect 17802 22820 17858 22822
rect 17562 21786 17618 21788
rect 17642 21786 17698 21788
rect 17722 21786 17778 21788
rect 17802 21786 17858 21788
rect 17562 21734 17588 21786
rect 17588 21734 17618 21786
rect 17642 21734 17652 21786
rect 17652 21734 17698 21786
rect 17722 21734 17768 21786
rect 17768 21734 17778 21786
rect 17802 21734 17832 21786
rect 17832 21734 17858 21786
rect 17562 21732 17618 21734
rect 17642 21732 17698 21734
rect 17722 21732 17778 21734
rect 17802 21732 17858 21734
rect 17562 20698 17618 20700
rect 17642 20698 17698 20700
rect 17722 20698 17778 20700
rect 17802 20698 17858 20700
rect 17562 20646 17588 20698
rect 17588 20646 17618 20698
rect 17642 20646 17652 20698
rect 17652 20646 17698 20698
rect 17722 20646 17768 20698
rect 17768 20646 17778 20698
rect 17802 20646 17832 20698
rect 17832 20646 17858 20698
rect 17562 20644 17618 20646
rect 17642 20644 17698 20646
rect 17722 20644 17778 20646
rect 17802 20644 17858 20646
rect 17562 19610 17618 19612
rect 17642 19610 17698 19612
rect 17722 19610 17778 19612
rect 17802 19610 17858 19612
rect 17562 19558 17588 19610
rect 17588 19558 17618 19610
rect 17642 19558 17652 19610
rect 17652 19558 17698 19610
rect 17722 19558 17768 19610
rect 17768 19558 17778 19610
rect 17802 19558 17832 19610
rect 17832 19558 17858 19610
rect 17562 19556 17618 19558
rect 17642 19556 17698 19558
rect 17722 19556 17778 19558
rect 17802 19556 17858 19558
rect 17314 19216 17370 19272
rect 16670 18536 16726 18592
rect 6491 2202 6547 2204
rect 6571 2202 6627 2204
rect 6651 2202 6707 2204
rect 6731 2202 6787 2204
rect 6491 2150 6517 2202
rect 6517 2150 6547 2202
rect 6571 2150 6581 2202
rect 6581 2150 6627 2202
rect 6651 2150 6697 2202
rect 6697 2150 6707 2202
rect 6731 2150 6761 2202
rect 6761 2150 6787 2202
rect 6491 2148 6547 2150
rect 6571 2148 6627 2150
rect 6651 2148 6707 2150
rect 6731 2148 6787 2150
rect 17562 18522 17618 18524
rect 17642 18522 17698 18524
rect 17722 18522 17778 18524
rect 17802 18522 17858 18524
rect 17562 18470 17588 18522
rect 17588 18470 17618 18522
rect 17642 18470 17652 18522
rect 17652 18470 17698 18522
rect 17722 18470 17768 18522
rect 17768 18470 17778 18522
rect 17802 18470 17832 18522
rect 17832 18470 17858 18522
rect 17562 18468 17618 18470
rect 17642 18468 17698 18470
rect 17722 18468 17778 18470
rect 17802 18468 17858 18470
rect 17562 17434 17618 17436
rect 17642 17434 17698 17436
rect 17722 17434 17778 17436
rect 17802 17434 17858 17436
rect 17562 17382 17588 17434
rect 17588 17382 17618 17434
rect 17642 17382 17652 17434
rect 17652 17382 17698 17434
rect 17722 17382 17768 17434
rect 17768 17382 17778 17434
rect 17802 17382 17832 17434
rect 17832 17382 17858 17434
rect 17562 17380 17618 17382
rect 17642 17380 17698 17382
rect 17722 17380 17778 17382
rect 17802 17380 17858 17382
rect 17562 16346 17618 16348
rect 17642 16346 17698 16348
rect 17722 16346 17778 16348
rect 17802 16346 17858 16348
rect 17562 16294 17588 16346
rect 17588 16294 17618 16346
rect 17642 16294 17652 16346
rect 17652 16294 17698 16346
rect 17722 16294 17768 16346
rect 17768 16294 17778 16346
rect 17802 16294 17832 16346
rect 17832 16294 17858 16346
rect 17562 16292 17618 16294
rect 17642 16292 17698 16294
rect 17722 16292 17778 16294
rect 17802 16292 17858 16294
rect 17562 15258 17618 15260
rect 17642 15258 17698 15260
rect 17722 15258 17778 15260
rect 17802 15258 17858 15260
rect 17562 15206 17588 15258
rect 17588 15206 17618 15258
rect 17642 15206 17652 15258
rect 17652 15206 17698 15258
rect 17722 15206 17768 15258
rect 17768 15206 17778 15258
rect 17802 15206 17832 15258
rect 17832 15206 17858 15258
rect 17562 15204 17618 15206
rect 17642 15204 17698 15206
rect 17722 15204 17778 15206
rect 17802 15204 17858 15206
rect 17562 14170 17618 14172
rect 17642 14170 17698 14172
rect 17722 14170 17778 14172
rect 17802 14170 17858 14172
rect 17562 14118 17588 14170
rect 17588 14118 17618 14170
rect 17642 14118 17652 14170
rect 17652 14118 17698 14170
rect 17722 14118 17768 14170
rect 17768 14118 17778 14170
rect 17802 14118 17832 14170
rect 17832 14118 17858 14170
rect 17562 14116 17618 14118
rect 17642 14116 17698 14118
rect 17722 14116 17778 14118
rect 17802 14116 17858 14118
rect 17562 13082 17618 13084
rect 17642 13082 17698 13084
rect 17722 13082 17778 13084
rect 17802 13082 17858 13084
rect 17562 13030 17588 13082
rect 17588 13030 17618 13082
rect 17642 13030 17652 13082
rect 17652 13030 17698 13082
rect 17722 13030 17768 13082
rect 17768 13030 17778 13082
rect 17802 13030 17832 13082
rect 17832 13030 17858 13082
rect 17562 13028 17618 13030
rect 17642 13028 17698 13030
rect 17722 13028 17778 13030
rect 17802 13028 17858 13030
rect 17562 11994 17618 11996
rect 17642 11994 17698 11996
rect 17722 11994 17778 11996
rect 17802 11994 17858 11996
rect 17562 11942 17588 11994
rect 17588 11942 17618 11994
rect 17642 11942 17652 11994
rect 17652 11942 17698 11994
rect 17722 11942 17768 11994
rect 17768 11942 17778 11994
rect 17802 11942 17832 11994
rect 17832 11942 17858 11994
rect 17562 11940 17618 11942
rect 17642 11940 17698 11942
rect 17722 11940 17778 11942
rect 17802 11940 17858 11942
rect 17562 10906 17618 10908
rect 17642 10906 17698 10908
rect 17722 10906 17778 10908
rect 17802 10906 17858 10908
rect 17562 10854 17588 10906
rect 17588 10854 17618 10906
rect 17642 10854 17652 10906
rect 17652 10854 17698 10906
rect 17722 10854 17768 10906
rect 17768 10854 17778 10906
rect 17802 10854 17832 10906
rect 17832 10854 17858 10906
rect 17562 10852 17618 10854
rect 17642 10852 17698 10854
rect 17722 10852 17778 10854
rect 17802 10852 17858 10854
rect 19890 18828 19946 18864
rect 19890 18808 19892 18828
rect 19892 18808 19944 18828
rect 19944 18808 19946 18828
rect 17562 9818 17618 9820
rect 17642 9818 17698 9820
rect 17722 9818 17778 9820
rect 17802 9818 17858 9820
rect 17562 9766 17588 9818
rect 17588 9766 17618 9818
rect 17642 9766 17652 9818
rect 17652 9766 17698 9818
rect 17722 9766 17768 9818
rect 17768 9766 17778 9818
rect 17802 9766 17832 9818
rect 17832 9766 17858 9818
rect 17562 9764 17618 9766
rect 17642 9764 17698 9766
rect 17722 9764 17778 9766
rect 17802 9764 17858 9766
rect 17562 8730 17618 8732
rect 17642 8730 17698 8732
rect 17722 8730 17778 8732
rect 17802 8730 17858 8732
rect 17562 8678 17588 8730
rect 17588 8678 17618 8730
rect 17642 8678 17652 8730
rect 17652 8678 17698 8730
rect 17722 8678 17768 8730
rect 17768 8678 17778 8730
rect 17802 8678 17832 8730
rect 17832 8678 17858 8730
rect 17562 8676 17618 8678
rect 17642 8676 17698 8678
rect 17722 8676 17778 8678
rect 17802 8676 17858 8678
rect 17562 7642 17618 7644
rect 17642 7642 17698 7644
rect 17722 7642 17778 7644
rect 17802 7642 17858 7644
rect 17562 7590 17588 7642
rect 17588 7590 17618 7642
rect 17642 7590 17652 7642
rect 17652 7590 17698 7642
rect 17722 7590 17768 7642
rect 17768 7590 17778 7642
rect 17802 7590 17832 7642
rect 17832 7590 17858 7642
rect 17562 7588 17618 7590
rect 17642 7588 17698 7590
rect 17722 7588 17778 7590
rect 17802 7588 17858 7590
rect 17562 6554 17618 6556
rect 17642 6554 17698 6556
rect 17722 6554 17778 6556
rect 17802 6554 17858 6556
rect 17562 6502 17588 6554
rect 17588 6502 17618 6554
rect 17642 6502 17652 6554
rect 17652 6502 17698 6554
rect 17722 6502 17768 6554
rect 17768 6502 17778 6554
rect 17802 6502 17832 6554
rect 17832 6502 17858 6554
rect 17562 6500 17618 6502
rect 17642 6500 17698 6502
rect 17722 6500 17778 6502
rect 17802 6500 17858 6502
rect 17562 5466 17618 5468
rect 17642 5466 17698 5468
rect 17722 5466 17778 5468
rect 17802 5466 17858 5468
rect 17562 5414 17588 5466
rect 17588 5414 17618 5466
rect 17642 5414 17652 5466
rect 17652 5414 17698 5466
rect 17722 5414 17768 5466
rect 17768 5414 17778 5466
rect 17802 5414 17832 5466
rect 17832 5414 17858 5466
rect 17562 5412 17618 5414
rect 17642 5412 17698 5414
rect 17722 5412 17778 5414
rect 17802 5412 17858 5414
rect 17562 4378 17618 4380
rect 17642 4378 17698 4380
rect 17722 4378 17778 4380
rect 17802 4378 17858 4380
rect 17562 4326 17588 4378
rect 17588 4326 17618 4378
rect 17642 4326 17652 4378
rect 17652 4326 17698 4378
rect 17722 4326 17768 4378
rect 17768 4326 17778 4378
rect 17802 4326 17832 4378
rect 17832 4326 17858 4378
rect 17562 4324 17618 4326
rect 17642 4324 17698 4326
rect 17722 4324 17778 4326
rect 17802 4324 17858 4326
rect 28632 34842 28688 34844
rect 28712 34842 28768 34844
rect 28792 34842 28848 34844
rect 28872 34842 28928 34844
rect 28632 34790 28658 34842
rect 28658 34790 28688 34842
rect 28712 34790 28722 34842
rect 28722 34790 28768 34842
rect 28792 34790 28838 34842
rect 28838 34790 28848 34842
rect 28872 34790 28902 34842
rect 28902 34790 28928 34842
rect 28632 34788 28688 34790
rect 28712 34788 28768 34790
rect 28792 34788 28848 34790
rect 28872 34788 28928 34790
rect 23097 34298 23153 34300
rect 23177 34298 23233 34300
rect 23257 34298 23313 34300
rect 23337 34298 23393 34300
rect 23097 34246 23123 34298
rect 23123 34246 23153 34298
rect 23177 34246 23187 34298
rect 23187 34246 23233 34298
rect 23257 34246 23303 34298
rect 23303 34246 23313 34298
rect 23337 34246 23367 34298
rect 23367 34246 23393 34298
rect 23097 34244 23153 34246
rect 23177 34244 23233 34246
rect 23257 34244 23313 34246
rect 23337 34244 23393 34246
rect 23097 33210 23153 33212
rect 23177 33210 23233 33212
rect 23257 33210 23313 33212
rect 23337 33210 23393 33212
rect 23097 33158 23123 33210
rect 23123 33158 23153 33210
rect 23177 33158 23187 33210
rect 23187 33158 23233 33210
rect 23257 33158 23303 33210
rect 23303 33158 23313 33210
rect 23337 33158 23367 33210
rect 23367 33158 23393 33210
rect 23097 33156 23153 33158
rect 23177 33156 23233 33158
rect 23257 33156 23313 33158
rect 23337 33156 23393 33158
rect 23097 32122 23153 32124
rect 23177 32122 23233 32124
rect 23257 32122 23313 32124
rect 23337 32122 23393 32124
rect 23097 32070 23123 32122
rect 23123 32070 23153 32122
rect 23177 32070 23187 32122
rect 23187 32070 23233 32122
rect 23257 32070 23303 32122
rect 23303 32070 23313 32122
rect 23337 32070 23367 32122
rect 23367 32070 23393 32122
rect 23097 32068 23153 32070
rect 23177 32068 23233 32070
rect 23257 32068 23313 32070
rect 23337 32068 23393 32070
rect 23097 31034 23153 31036
rect 23177 31034 23233 31036
rect 23257 31034 23313 31036
rect 23337 31034 23393 31036
rect 23097 30982 23123 31034
rect 23123 30982 23153 31034
rect 23177 30982 23187 31034
rect 23187 30982 23233 31034
rect 23257 30982 23303 31034
rect 23303 30982 23313 31034
rect 23337 30982 23367 31034
rect 23367 30982 23393 31034
rect 23097 30980 23153 30982
rect 23177 30980 23233 30982
rect 23257 30980 23313 30982
rect 23337 30980 23393 30982
rect 28632 33754 28688 33756
rect 28712 33754 28768 33756
rect 28792 33754 28848 33756
rect 28872 33754 28928 33756
rect 28632 33702 28658 33754
rect 28658 33702 28688 33754
rect 28712 33702 28722 33754
rect 28722 33702 28768 33754
rect 28792 33702 28838 33754
rect 28838 33702 28848 33754
rect 28872 33702 28902 33754
rect 28902 33702 28928 33754
rect 28632 33700 28688 33702
rect 28712 33700 28768 33702
rect 28792 33700 28848 33702
rect 28872 33700 28928 33702
rect 23097 29946 23153 29948
rect 23177 29946 23233 29948
rect 23257 29946 23313 29948
rect 23337 29946 23393 29948
rect 23097 29894 23123 29946
rect 23123 29894 23153 29946
rect 23177 29894 23187 29946
rect 23187 29894 23233 29946
rect 23257 29894 23303 29946
rect 23303 29894 23313 29946
rect 23337 29894 23367 29946
rect 23367 29894 23393 29946
rect 23097 29892 23153 29894
rect 23177 29892 23233 29894
rect 23257 29892 23313 29894
rect 23337 29892 23393 29894
rect 23097 28858 23153 28860
rect 23177 28858 23233 28860
rect 23257 28858 23313 28860
rect 23337 28858 23393 28860
rect 23097 28806 23123 28858
rect 23123 28806 23153 28858
rect 23177 28806 23187 28858
rect 23187 28806 23233 28858
rect 23257 28806 23303 28858
rect 23303 28806 23313 28858
rect 23337 28806 23367 28858
rect 23367 28806 23393 28858
rect 23097 28804 23153 28806
rect 23177 28804 23233 28806
rect 23257 28804 23313 28806
rect 23337 28804 23393 28806
rect 20626 19372 20682 19408
rect 20626 19352 20628 19372
rect 20628 19352 20680 19372
rect 20680 19352 20682 19372
rect 23097 27770 23153 27772
rect 23177 27770 23233 27772
rect 23257 27770 23313 27772
rect 23337 27770 23393 27772
rect 23097 27718 23123 27770
rect 23123 27718 23153 27770
rect 23177 27718 23187 27770
rect 23187 27718 23233 27770
rect 23257 27718 23303 27770
rect 23303 27718 23313 27770
rect 23337 27718 23367 27770
rect 23367 27718 23393 27770
rect 23097 27716 23153 27718
rect 23177 27716 23233 27718
rect 23257 27716 23313 27718
rect 23337 27716 23393 27718
rect 23097 26682 23153 26684
rect 23177 26682 23233 26684
rect 23257 26682 23313 26684
rect 23337 26682 23393 26684
rect 23097 26630 23123 26682
rect 23123 26630 23153 26682
rect 23177 26630 23187 26682
rect 23187 26630 23233 26682
rect 23257 26630 23303 26682
rect 23303 26630 23313 26682
rect 23337 26630 23367 26682
rect 23367 26630 23393 26682
rect 23097 26628 23153 26630
rect 23177 26628 23233 26630
rect 23257 26628 23313 26630
rect 23337 26628 23393 26630
rect 23097 25594 23153 25596
rect 23177 25594 23233 25596
rect 23257 25594 23313 25596
rect 23337 25594 23393 25596
rect 23097 25542 23123 25594
rect 23123 25542 23153 25594
rect 23177 25542 23187 25594
rect 23187 25542 23233 25594
rect 23257 25542 23303 25594
rect 23303 25542 23313 25594
rect 23337 25542 23367 25594
rect 23367 25542 23393 25594
rect 23097 25540 23153 25542
rect 23177 25540 23233 25542
rect 23257 25540 23313 25542
rect 23337 25540 23393 25542
rect 23097 24506 23153 24508
rect 23177 24506 23233 24508
rect 23257 24506 23313 24508
rect 23337 24506 23393 24508
rect 23097 24454 23123 24506
rect 23123 24454 23153 24506
rect 23177 24454 23187 24506
rect 23187 24454 23233 24506
rect 23257 24454 23303 24506
rect 23303 24454 23313 24506
rect 23337 24454 23367 24506
rect 23367 24454 23393 24506
rect 23097 24452 23153 24454
rect 23177 24452 23233 24454
rect 23257 24452 23313 24454
rect 23337 24452 23393 24454
rect 23097 23418 23153 23420
rect 23177 23418 23233 23420
rect 23257 23418 23313 23420
rect 23337 23418 23393 23420
rect 23097 23366 23123 23418
rect 23123 23366 23153 23418
rect 23177 23366 23187 23418
rect 23187 23366 23233 23418
rect 23257 23366 23303 23418
rect 23303 23366 23313 23418
rect 23337 23366 23367 23418
rect 23367 23366 23393 23418
rect 23097 23364 23153 23366
rect 23177 23364 23233 23366
rect 23257 23364 23313 23366
rect 23337 23364 23393 23366
rect 23097 22330 23153 22332
rect 23177 22330 23233 22332
rect 23257 22330 23313 22332
rect 23337 22330 23393 22332
rect 23097 22278 23123 22330
rect 23123 22278 23153 22330
rect 23177 22278 23187 22330
rect 23187 22278 23233 22330
rect 23257 22278 23303 22330
rect 23303 22278 23313 22330
rect 23337 22278 23367 22330
rect 23367 22278 23393 22330
rect 23097 22276 23153 22278
rect 23177 22276 23233 22278
rect 23257 22276 23313 22278
rect 23337 22276 23393 22278
rect 22466 19372 22522 19408
rect 22466 19352 22468 19372
rect 22468 19352 22520 19372
rect 22520 19352 22522 19372
rect 23097 21242 23153 21244
rect 23177 21242 23233 21244
rect 23257 21242 23313 21244
rect 23337 21242 23393 21244
rect 23097 21190 23123 21242
rect 23123 21190 23153 21242
rect 23177 21190 23187 21242
rect 23187 21190 23233 21242
rect 23257 21190 23303 21242
rect 23303 21190 23313 21242
rect 23337 21190 23367 21242
rect 23367 21190 23393 21242
rect 23097 21188 23153 21190
rect 23177 21188 23233 21190
rect 23257 21188 23313 21190
rect 23337 21188 23393 21190
rect 23097 20154 23153 20156
rect 23177 20154 23233 20156
rect 23257 20154 23313 20156
rect 23337 20154 23393 20156
rect 23097 20102 23123 20154
rect 23123 20102 23153 20154
rect 23177 20102 23187 20154
rect 23187 20102 23233 20154
rect 23257 20102 23303 20154
rect 23303 20102 23313 20154
rect 23337 20102 23367 20154
rect 23367 20102 23393 20154
rect 23097 20100 23153 20102
rect 23177 20100 23233 20102
rect 23257 20100 23313 20102
rect 23337 20100 23393 20102
rect 17562 3290 17618 3292
rect 17642 3290 17698 3292
rect 17722 3290 17778 3292
rect 17802 3290 17858 3292
rect 17562 3238 17588 3290
rect 17588 3238 17618 3290
rect 17642 3238 17652 3290
rect 17652 3238 17698 3290
rect 17722 3238 17768 3290
rect 17768 3238 17778 3290
rect 17802 3238 17832 3290
rect 17832 3238 17858 3290
rect 17562 3236 17618 3238
rect 17642 3236 17698 3238
rect 17722 3236 17778 3238
rect 17802 3236 17858 3238
rect 23097 19066 23153 19068
rect 23177 19066 23233 19068
rect 23257 19066 23313 19068
rect 23337 19066 23393 19068
rect 23097 19014 23123 19066
rect 23123 19014 23153 19066
rect 23177 19014 23187 19066
rect 23187 19014 23233 19066
rect 23257 19014 23303 19066
rect 23303 19014 23313 19066
rect 23337 19014 23367 19066
rect 23367 19014 23393 19066
rect 23097 19012 23153 19014
rect 23177 19012 23233 19014
rect 23257 19012 23313 19014
rect 23337 19012 23393 19014
rect 23097 17978 23153 17980
rect 23177 17978 23233 17980
rect 23257 17978 23313 17980
rect 23337 17978 23393 17980
rect 23097 17926 23123 17978
rect 23123 17926 23153 17978
rect 23177 17926 23187 17978
rect 23187 17926 23233 17978
rect 23257 17926 23303 17978
rect 23303 17926 23313 17978
rect 23337 17926 23367 17978
rect 23367 17926 23393 17978
rect 23097 17924 23153 17926
rect 23177 17924 23233 17926
rect 23257 17924 23313 17926
rect 23337 17924 23393 17926
rect 23097 16890 23153 16892
rect 23177 16890 23233 16892
rect 23257 16890 23313 16892
rect 23337 16890 23393 16892
rect 23097 16838 23123 16890
rect 23123 16838 23153 16890
rect 23177 16838 23187 16890
rect 23187 16838 23233 16890
rect 23257 16838 23303 16890
rect 23303 16838 23313 16890
rect 23337 16838 23367 16890
rect 23367 16838 23393 16890
rect 23097 16836 23153 16838
rect 23177 16836 23233 16838
rect 23257 16836 23313 16838
rect 23337 16836 23393 16838
rect 28632 32666 28688 32668
rect 28712 32666 28768 32668
rect 28792 32666 28848 32668
rect 28872 32666 28928 32668
rect 28632 32614 28658 32666
rect 28658 32614 28688 32666
rect 28712 32614 28722 32666
rect 28722 32614 28768 32666
rect 28792 32614 28838 32666
rect 28838 32614 28848 32666
rect 28872 32614 28902 32666
rect 28902 32614 28928 32666
rect 28632 32612 28688 32614
rect 28712 32612 28768 32614
rect 28792 32612 28848 32614
rect 28872 32612 28928 32614
rect 25594 18808 25650 18864
rect 23097 15802 23153 15804
rect 23177 15802 23233 15804
rect 23257 15802 23313 15804
rect 23337 15802 23393 15804
rect 23097 15750 23123 15802
rect 23123 15750 23153 15802
rect 23177 15750 23187 15802
rect 23187 15750 23233 15802
rect 23257 15750 23303 15802
rect 23303 15750 23313 15802
rect 23337 15750 23367 15802
rect 23367 15750 23393 15802
rect 23097 15748 23153 15750
rect 23177 15748 23233 15750
rect 23257 15748 23313 15750
rect 23337 15748 23393 15750
rect 23097 14714 23153 14716
rect 23177 14714 23233 14716
rect 23257 14714 23313 14716
rect 23337 14714 23393 14716
rect 23097 14662 23123 14714
rect 23123 14662 23153 14714
rect 23177 14662 23187 14714
rect 23187 14662 23233 14714
rect 23257 14662 23303 14714
rect 23303 14662 23313 14714
rect 23337 14662 23367 14714
rect 23367 14662 23393 14714
rect 23097 14660 23153 14662
rect 23177 14660 23233 14662
rect 23257 14660 23313 14662
rect 23337 14660 23393 14662
rect 23097 13626 23153 13628
rect 23177 13626 23233 13628
rect 23257 13626 23313 13628
rect 23337 13626 23393 13628
rect 23097 13574 23123 13626
rect 23123 13574 23153 13626
rect 23177 13574 23187 13626
rect 23187 13574 23233 13626
rect 23257 13574 23303 13626
rect 23303 13574 23313 13626
rect 23337 13574 23367 13626
rect 23367 13574 23393 13626
rect 23097 13572 23153 13574
rect 23177 13572 23233 13574
rect 23257 13572 23313 13574
rect 23337 13572 23393 13574
rect 23097 12538 23153 12540
rect 23177 12538 23233 12540
rect 23257 12538 23313 12540
rect 23337 12538 23393 12540
rect 23097 12486 23123 12538
rect 23123 12486 23153 12538
rect 23177 12486 23187 12538
rect 23187 12486 23233 12538
rect 23257 12486 23303 12538
rect 23303 12486 23313 12538
rect 23337 12486 23367 12538
rect 23367 12486 23393 12538
rect 23097 12484 23153 12486
rect 23177 12484 23233 12486
rect 23257 12484 23313 12486
rect 23337 12484 23393 12486
rect 23097 11450 23153 11452
rect 23177 11450 23233 11452
rect 23257 11450 23313 11452
rect 23337 11450 23393 11452
rect 23097 11398 23123 11450
rect 23123 11398 23153 11450
rect 23177 11398 23187 11450
rect 23187 11398 23233 11450
rect 23257 11398 23303 11450
rect 23303 11398 23313 11450
rect 23337 11398 23367 11450
rect 23367 11398 23393 11450
rect 23097 11396 23153 11398
rect 23177 11396 23233 11398
rect 23257 11396 23313 11398
rect 23337 11396 23393 11398
rect 23097 10362 23153 10364
rect 23177 10362 23233 10364
rect 23257 10362 23313 10364
rect 23337 10362 23393 10364
rect 23097 10310 23123 10362
rect 23123 10310 23153 10362
rect 23177 10310 23187 10362
rect 23187 10310 23233 10362
rect 23257 10310 23303 10362
rect 23303 10310 23313 10362
rect 23337 10310 23367 10362
rect 23367 10310 23393 10362
rect 23097 10308 23153 10310
rect 23177 10308 23233 10310
rect 23257 10308 23313 10310
rect 23337 10308 23393 10310
rect 23097 9274 23153 9276
rect 23177 9274 23233 9276
rect 23257 9274 23313 9276
rect 23337 9274 23393 9276
rect 23097 9222 23123 9274
rect 23123 9222 23153 9274
rect 23177 9222 23187 9274
rect 23187 9222 23233 9274
rect 23257 9222 23303 9274
rect 23303 9222 23313 9274
rect 23337 9222 23367 9274
rect 23367 9222 23393 9274
rect 23097 9220 23153 9222
rect 23177 9220 23233 9222
rect 23257 9220 23313 9222
rect 23337 9220 23393 9222
rect 23097 8186 23153 8188
rect 23177 8186 23233 8188
rect 23257 8186 23313 8188
rect 23337 8186 23393 8188
rect 23097 8134 23123 8186
rect 23123 8134 23153 8186
rect 23177 8134 23187 8186
rect 23187 8134 23233 8186
rect 23257 8134 23303 8186
rect 23303 8134 23313 8186
rect 23337 8134 23367 8186
rect 23367 8134 23393 8186
rect 23097 8132 23153 8134
rect 23177 8132 23233 8134
rect 23257 8132 23313 8134
rect 23337 8132 23393 8134
rect 23097 7098 23153 7100
rect 23177 7098 23233 7100
rect 23257 7098 23313 7100
rect 23337 7098 23393 7100
rect 23097 7046 23123 7098
rect 23123 7046 23153 7098
rect 23177 7046 23187 7098
rect 23187 7046 23233 7098
rect 23257 7046 23303 7098
rect 23303 7046 23313 7098
rect 23337 7046 23367 7098
rect 23367 7046 23393 7098
rect 23097 7044 23153 7046
rect 23177 7044 23233 7046
rect 23257 7044 23313 7046
rect 23337 7044 23393 7046
rect 23097 6010 23153 6012
rect 23177 6010 23233 6012
rect 23257 6010 23313 6012
rect 23337 6010 23393 6012
rect 23097 5958 23123 6010
rect 23123 5958 23153 6010
rect 23177 5958 23187 6010
rect 23187 5958 23233 6010
rect 23257 5958 23303 6010
rect 23303 5958 23313 6010
rect 23337 5958 23367 6010
rect 23367 5958 23393 6010
rect 23097 5956 23153 5958
rect 23177 5956 23233 5958
rect 23257 5956 23313 5958
rect 23337 5956 23393 5958
rect 23097 4922 23153 4924
rect 23177 4922 23233 4924
rect 23257 4922 23313 4924
rect 23337 4922 23393 4924
rect 23097 4870 23123 4922
rect 23123 4870 23153 4922
rect 23177 4870 23187 4922
rect 23187 4870 23233 4922
rect 23257 4870 23303 4922
rect 23303 4870 23313 4922
rect 23337 4870 23367 4922
rect 23367 4870 23393 4922
rect 23097 4868 23153 4870
rect 23177 4868 23233 4870
rect 23257 4868 23313 4870
rect 23337 4868 23393 4870
rect 23097 3834 23153 3836
rect 23177 3834 23233 3836
rect 23257 3834 23313 3836
rect 23337 3834 23393 3836
rect 23097 3782 23123 3834
rect 23123 3782 23153 3834
rect 23177 3782 23187 3834
rect 23187 3782 23233 3834
rect 23257 3782 23303 3834
rect 23303 3782 23313 3834
rect 23337 3782 23367 3834
rect 23367 3782 23393 3834
rect 23097 3780 23153 3782
rect 23177 3780 23233 3782
rect 23257 3780 23313 3782
rect 23337 3780 23393 3782
rect 28632 31578 28688 31580
rect 28712 31578 28768 31580
rect 28792 31578 28848 31580
rect 28872 31578 28928 31580
rect 28632 31526 28658 31578
rect 28658 31526 28688 31578
rect 28712 31526 28722 31578
rect 28722 31526 28768 31578
rect 28792 31526 28838 31578
rect 28838 31526 28848 31578
rect 28872 31526 28902 31578
rect 28902 31526 28928 31578
rect 28632 31524 28688 31526
rect 28712 31524 28768 31526
rect 28792 31524 28848 31526
rect 28872 31524 28928 31526
rect 28632 30490 28688 30492
rect 28712 30490 28768 30492
rect 28792 30490 28848 30492
rect 28872 30490 28928 30492
rect 28632 30438 28658 30490
rect 28658 30438 28688 30490
rect 28712 30438 28722 30490
rect 28722 30438 28768 30490
rect 28792 30438 28838 30490
rect 28838 30438 28848 30490
rect 28872 30438 28902 30490
rect 28902 30438 28928 30490
rect 28632 30436 28688 30438
rect 28712 30436 28768 30438
rect 28792 30436 28848 30438
rect 28872 30436 28928 30438
rect 28632 29402 28688 29404
rect 28712 29402 28768 29404
rect 28792 29402 28848 29404
rect 28872 29402 28928 29404
rect 28632 29350 28658 29402
rect 28658 29350 28688 29402
rect 28712 29350 28722 29402
rect 28722 29350 28768 29402
rect 28792 29350 28838 29402
rect 28838 29350 28848 29402
rect 28872 29350 28902 29402
rect 28902 29350 28928 29402
rect 28632 29348 28688 29350
rect 28712 29348 28768 29350
rect 28792 29348 28848 29350
rect 28872 29348 28928 29350
rect 28632 28314 28688 28316
rect 28712 28314 28768 28316
rect 28792 28314 28848 28316
rect 28872 28314 28928 28316
rect 28632 28262 28658 28314
rect 28658 28262 28688 28314
rect 28712 28262 28722 28314
rect 28722 28262 28768 28314
rect 28792 28262 28838 28314
rect 28838 28262 28848 28314
rect 28872 28262 28902 28314
rect 28902 28262 28928 28314
rect 28632 28260 28688 28262
rect 28712 28260 28768 28262
rect 28792 28260 28848 28262
rect 28872 28260 28928 28262
rect 28632 27226 28688 27228
rect 28712 27226 28768 27228
rect 28792 27226 28848 27228
rect 28872 27226 28928 27228
rect 28632 27174 28658 27226
rect 28658 27174 28688 27226
rect 28712 27174 28722 27226
rect 28722 27174 28768 27226
rect 28792 27174 28838 27226
rect 28838 27174 28848 27226
rect 28872 27174 28902 27226
rect 28902 27174 28928 27226
rect 28632 27172 28688 27174
rect 28712 27172 28768 27174
rect 28792 27172 28848 27174
rect 28872 27172 28928 27174
rect 28632 26138 28688 26140
rect 28712 26138 28768 26140
rect 28792 26138 28848 26140
rect 28872 26138 28928 26140
rect 28632 26086 28658 26138
rect 28658 26086 28688 26138
rect 28712 26086 28722 26138
rect 28722 26086 28768 26138
rect 28792 26086 28838 26138
rect 28838 26086 28848 26138
rect 28872 26086 28902 26138
rect 28902 26086 28928 26138
rect 28632 26084 28688 26086
rect 28712 26084 28768 26086
rect 28792 26084 28848 26086
rect 28872 26084 28928 26086
rect 28632 25050 28688 25052
rect 28712 25050 28768 25052
rect 28792 25050 28848 25052
rect 28872 25050 28928 25052
rect 28632 24998 28658 25050
rect 28658 24998 28688 25050
rect 28712 24998 28722 25050
rect 28722 24998 28768 25050
rect 28792 24998 28838 25050
rect 28838 24998 28848 25050
rect 28872 24998 28902 25050
rect 28902 24998 28928 25050
rect 28632 24996 28688 24998
rect 28712 24996 28768 24998
rect 28792 24996 28848 24998
rect 28872 24996 28928 24998
rect 28632 23962 28688 23964
rect 28712 23962 28768 23964
rect 28792 23962 28848 23964
rect 28872 23962 28928 23964
rect 28632 23910 28658 23962
rect 28658 23910 28688 23962
rect 28712 23910 28722 23962
rect 28722 23910 28768 23962
rect 28792 23910 28838 23962
rect 28838 23910 28848 23962
rect 28872 23910 28902 23962
rect 28902 23910 28928 23962
rect 28632 23908 28688 23910
rect 28712 23908 28768 23910
rect 28792 23908 28848 23910
rect 28872 23908 28928 23910
rect 28632 22874 28688 22876
rect 28712 22874 28768 22876
rect 28792 22874 28848 22876
rect 28872 22874 28928 22876
rect 28632 22822 28658 22874
rect 28658 22822 28688 22874
rect 28712 22822 28722 22874
rect 28722 22822 28768 22874
rect 28792 22822 28838 22874
rect 28838 22822 28848 22874
rect 28872 22822 28902 22874
rect 28902 22822 28928 22874
rect 28632 22820 28688 22822
rect 28712 22820 28768 22822
rect 28792 22820 28848 22822
rect 28872 22820 28928 22822
rect 28632 21786 28688 21788
rect 28712 21786 28768 21788
rect 28792 21786 28848 21788
rect 28872 21786 28928 21788
rect 28632 21734 28658 21786
rect 28658 21734 28688 21786
rect 28712 21734 28722 21786
rect 28722 21734 28768 21786
rect 28792 21734 28838 21786
rect 28838 21734 28848 21786
rect 28872 21734 28902 21786
rect 28902 21734 28928 21786
rect 28632 21732 28688 21734
rect 28712 21732 28768 21734
rect 28792 21732 28848 21734
rect 28872 21732 28928 21734
rect 28632 20698 28688 20700
rect 28712 20698 28768 20700
rect 28792 20698 28848 20700
rect 28872 20698 28928 20700
rect 28632 20646 28658 20698
rect 28658 20646 28688 20698
rect 28712 20646 28722 20698
rect 28722 20646 28768 20698
rect 28792 20646 28838 20698
rect 28838 20646 28848 20698
rect 28872 20646 28902 20698
rect 28902 20646 28928 20698
rect 28632 20644 28688 20646
rect 28712 20644 28768 20646
rect 28792 20644 28848 20646
rect 28872 20644 28928 20646
rect 28632 19610 28688 19612
rect 28712 19610 28768 19612
rect 28792 19610 28848 19612
rect 28872 19610 28928 19612
rect 28632 19558 28658 19610
rect 28658 19558 28688 19610
rect 28712 19558 28722 19610
rect 28722 19558 28768 19610
rect 28792 19558 28838 19610
rect 28838 19558 28848 19610
rect 28872 19558 28902 19610
rect 28902 19558 28928 19610
rect 28632 19556 28688 19558
rect 28712 19556 28768 19558
rect 28792 19556 28848 19558
rect 28872 19556 28928 19558
rect 28632 18522 28688 18524
rect 28712 18522 28768 18524
rect 28792 18522 28848 18524
rect 28872 18522 28928 18524
rect 28632 18470 28658 18522
rect 28658 18470 28688 18522
rect 28712 18470 28722 18522
rect 28722 18470 28768 18522
rect 28792 18470 28838 18522
rect 28838 18470 28848 18522
rect 28872 18470 28902 18522
rect 28902 18470 28928 18522
rect 28632 18468 28688 18470
rect 28712 18468 28768 18470
rect 28792 18468 28848 18470
rect 28872 18468 28928 18470
rect 28632 17434 28688 17436
rect 28712 17434 28768 17436
rect 28792 17434 28848 17436
rect 28872 17434 28928 17436
rect 28632 17382 28658 17434
rect 28658 17382 28688 17434
rect 28712 17382 28722 17434
rect 28722 17382 28768 17434
rect 28792 17382 28838 17434
rect 28838 17382 28848 17434
rect 28872 17382 28902 17434
rect 28902 17382 28928 17434
rect 28632 17380 28688 17382
rect 28712 17380 28768 17382
rect 28792 17380 28848 17382
rect 28872 17380 28928 17382
rect 28632 16346 28688 16348
rect 28712 16346 28768 16348
rect 28792 16346 28848 16348
rect 28872 16346 28928 16348
rect 28632 16294 28658 16346
rect 28658 16294 28688 16346
rect 28712 16294 28722 16346
rect 28722 16294 28768 16346
rect 28792 16294 28838 16346
rect 28838 16294 28848 16346
rect 28872 16294 28902 16346
rect 28902 16294 28928 16346
rect 28632 16292 28688 16294
rect 28712 16292 28768 16294
rect 28792 16292 28848 16294
rect 28872 16292 28928 16294
rect 28632 15258 28688 15260
rect 28712 15258 28768 15260
rect 28792 15258 28848 15260
rect 28872 15258 28928 15260
rect 28632 15206 28658 15258
rect 28658 15206 28688 15258
rect 28712 15206 28722 15258
rect 28722 15206 28768 15258
rect 28792 15206 28838 15258
rect 28838 15206 28848 15258
rect 28872 15206 28902 15258
rect 28902 15206 28928 15258
rect 28632 15204 28688 15206
rect 28712 15204 28768 15206
rect 28792 15204 28848 15206
rect 28872 15204 28928 15206
rect 28632 14170 28688 14172
rect 28712 14170 28768 14172
rect 28792 14170 28848 14172
rect 28872 14170 28928 14172
rect 28632 14118 28658 14170
rect 28658 14118 28688 14170
rect 28712 14118 28722 14170
rect 28722 14118 28768 14170
rect 28792 14118 28838 14170
rect 28838 14118 28848 14170
rect 28872 14118 28902 14170
rect 28902 14118 28928 14170
rect 28632 14116 28688 14118
rect 28712 14116 28768 14118
rect 28792 14116 28848 14118
rect 28872 14116 28928 14118
rect 28632 13082 28688 13084
rect 28712 13082 28768 13084
rect 28792 13082 28848 13084
rect 28872 13082 28928 13084
rect 28632 13030 28658 13082
rect 28658 13030 28688 13082
rect 28712 13030 28722 13082
rect 28722 13030 28768 13082
rect 28792 13030 28838 13082
rect 28838 13030 28848 13082
rect 28872 13030 28902 13082
rect 28902 13030 28928 13082
rect 28632 13028 28688 13030
rect 28712 13028 28768 13030
rect 28792 13028 28848 13030
rect 28872 13028 28928 13030
rect 28632 11994 28688 11996
rect 28712 11994 28768 11996
rect 28792 11994 28848 11996
rect 28872 11994 28928 11996
rect 28632 11942 28658 11994
rect 28658 11942 28688 11994
rect 28712 11942 28722 11994
rect 28722 11942 28768 11994
rect 28792 11942 28838 11994
rect 28838 11942 28848 11994
rect 28872 11942 28902 11994
rect 28902 11942 28928 11994
rect 28632 11940 28688 11942
rect 28712 11940 28768 11942
rect 28792 11940 28848 11942
rect 28872 11940 28928 11942
rect 28632 10906 28688 10908
rect 28712 10906 28768 10908
rect 28792 10906 28848 10908
rect 28872 10906 28928 10908
rect 28632 10854 28658 10906
rect 28658 10854 28688 10906
rect 28712 10854 28722 10906
rect 28722 10854 28768 10906
rect 28792 10854 28838 10906
rect 28838 10854 28848 10906
rect 28872 10854 28902 10906
rect 28902 10854 28928 10906
rect 28632 10852 28688 10854
rect 28712 10852 28768 10854
rect 28792 10852 28848 10854
rect 28872 10852 28928 10854
rect 28632 9818 28688 9820
rect 28712 9818 28768 9820
rect 28792 9818 28848 9820
rect 28872 9818 28928 9820
rect 28632 9766 28658 9818
rect 28658 9766 28688 9818
rect 28712 9766 28722 9818
rect 28722 9766 28768 9818
rect 28792 9766 28838 9818
rect 28838 9766 28848 9818
rect 28872 9766 28902 9818
rect 28902 9766 28928 9818
rect 28632 9764 28688 9766
rect 28712 9764 28768 9766
rect 28792 9764 28848 9766
rect 28872 9764 28928 9766
rect 28632 8730 28688 8732
rect 28712 8730 28768 8732
rect 28792 8730 28848 8732
rect 28872 8730 28928 8732
rect 28632 8678 28658 8730
rect 28658 8678 28688 8730
rect 28712 8678 28722 8730
rect 28722 8678 28768 8730
rect 28792 8678 28838 8730
rect 28838 8678 28848 8730
rect 28872 8678 28902 8730
rect 28902 8678 28928 8730
rect 28632 8676 28688 8678
rect 28712 8676 28768 8678
rect 28792 8676 28848 8678
rect 28872 8676 28928 8678
rect 28632 7642 28688 7644
rect 28712 7642 28768 7644
rect 28792 7642 28848 7644
rect 28872 7642 28928 7644
rect 28632 7590 28658 7642
rect 28658 7590 28688 7642
rect 28712 7590 28722 7642
rect 28722 7590 28768 7642
rect 28792 7590 28838 7642
rect 28838 7590 28848 7642
rect 28872 7590 28902 7642
rect 28902 7590 28928 7642
rect 28632 7588 28688 7590
rect 28712 7588 28768 7590
rect 28792 7588 28848 7590
rect 28872 7588 28928 7590
rect 28632 6554 28688 6556
rect 28712 6554 28768 6556
rect 28792 6554 28848 6556
rect 28872 6554 28928 6556
rect 28632 6502 28658 6554
rect 28658 6502 28688 6554
rect 28712 6502 28722 6554
rect 28722 6502 28768 6554
rect 28792 6502 28838 6554
rect 28838 6502 28848 6554
rect 28872 6502 28902 6554
rect 28902 6502 28928 6554
rect 28632 6500 28688 6502
rect 28712 6500 28768 6502
rect 28792 6500 28848 6502
rect 28872 6500 28928 6502
rect 30470 8880 30526 8936
rect 28632 5466 28688 5468
rect 28712 5466 28768 5468
rect 28792 5466 28848 5468
rect 28872 5466 28928 5468
rect 28632 5414 28658 5466
rect 28658 5414 28688 5466
rect 28712 5414 28722 5466
rect 28722 5414 28768 5466
rect 28792 5414 28838 5466
rect 28838 5414 28848 5466
rect 28872 5414 28902 5466
rect 28902 5414 28928 5466
rect 28632 5412 28688 5414
rect 28712 5412 28768 5414
rect 28792 5412 28848 5414
rect 28872 5412 28928 5414
rect 28632 4378 28688 4380
rect 28712 4378 28768 4380
rect 28792 4378 28848 4380
rect 28872 4378 28928 4380
rect 28632 4326 28658 4378
rect 28658 4326 28688 4378
rect 28712 4326 28722 4378
rect 28722 4326 28768 4378
rect 28792 4326 28838 4378
rect 28838 4326 28848 4378
rect 28872 4326 28902 4378
rect 28902 4326 28928 4378
rect 28632 4324 28688 4326
rect 28712 4324 28768 4326
rect 28792 4324 28848 4326
rect 28872 4324 28928 4326
rect 33598 33396 33600 33416
rect 33600 33396 33652 33416
rect 33652 33396 33654 33416
rect 33598 33360 33654 33396
rect 33598 29280 33654 29336
rect 33506 25200 33562 25256
rect 33598 21120 33654 21176
rect 33598 17060 33654 17096
rect 33598 17040 33600 17060
rect 33600 17040 33652 17060
rect 33652 17040 33654 17060
rect 33598 12960 33654 13016
rect 23097 2746 23153 2748
rect 23177 2746 23233 2748
rect 23257 2746 23313 2748
rect 23337 2746 23393 2748
rect 23097 2694 23123 2746
rect 23123 2694 23153 2746
rect 23177 2694 23187 2746
rect 23187 2694 23233 2746
rect 23257 2694 23303 2746
rect 23303 2694 23313 2746
rect 23337 2694 23367 2746
rect 23367 2694 23393 2746
rect 23097 2692 23153 2694
rect 23177 2692 23233 2694
rect 23257 2692 23313 2694
rect 23337 2692 23393 2694
rect 28632 3290 28688 3292
rect 28712 3290 28768 3292
rect 28792 3290 28848 3292
rect 28872 3290 28928 3292
rect 28632 3238 28658 3290
rect 28658 3238 28688 3290
rect 28712 3238 28722 3290
rect 28722 3238 28768 3290
rect 28792 3238 28838 3290
rect 28838 3238 28848 3290
rect 28872 3238 28902 3290
rect 28902 3238 28928 3290
rect 28632 3236 28688 3238
rect 28712 3236 28768 3238
rect 28792 3236 28848 3238
rect 28872 3236 28928 3238
rect 33598 4800 33654 4856
rect 17562 2202 17618 2204
rect 17642 2202 17698 2204
rect 17722 2202 17778 2204
rect 17802 2202 17858 2204
rect 17562 2150 17588 2202
rect 17588 2150 17618 2202
rect 17642 2150 17652 2202
rect 17652 2150 17698 2202
rect 17722 2150 17768 2202
rect 17768 2150 17778 2202
rect 17802 2150 17832 2202
rect 17832 2150 17858 2202
rect 17562 2148 17618 2150
rect 17642 2148 17698 2150
rect 17722 2148 17778 2150
rect 17802 2148 17858 2150
rect 28632 2202 28688 2204
rect 28712 2202 28768 2204
rect 28792 2202 28848 2204
rect 28872 2202 28928 2204
rect 28632 2150 28658 2202
rect 28658 2150 28688 2202
rect 28712 2150 28722 2202
rect 28722 2150 28768 2202
rect 28792 2150 28838 2202
rect 28838 2150 28848 2202
rect 28872 2150 28902 2202
rect 28902 2150 28928 2202
rect 28632 2148 28688 2150
rect 28712 2148 28768 2150
rect 28792 2148 28848 2150
rect 28872 2148 28928 2150
rect 31942 720 31998 776
<< metal3 >>
rect 0 36818 800 36848
rect 1393 36818 1459 36821
rect 0 36816 1459 36818
rect 0 36760 1398 36816
rect 1454 36760 1459 36816
rect 0 36758 1459 36760
rect 0 36728 800 36758
rect 1393 36755 1459 36758
rect 12014 35392 12334 35393
rect 12014 35328 12022 35392
rect 12086 35328 12102 35392
rect 12166 35328 12182 35392
rect 12246 35328 12262 35392
rect 12326 35328 12334 35392
rect 12014 35327 12334 35328
rect 23085 35392 23405 35393
rect 23085 35328 23093 35392
rect 23157 35328 23173 35392
rect 23237 35328 23253 35392
rect 23317 35328 23333 35392
rect 23397 35328 23405 35392
rect 23085 35327 23405 35328
rect 6479 34848 6799 34849
rect 6479 34784 6487 34848
rect 6551 34784 6567 34848
rect 6631 34784 6647 34848
rect 6711 34784 6727 34848
rect 6791 34784 6799 34848
rect 6479 34783 6799 34784
rect 17550 34848 17870 34849
rect 17550 34784 17558 34848
rect 17622 34784 17638 34848
rect 17702 34784 17718 34848
rect 17782 34784 17798 34848
rect 17862 34784 17870 34848
rect 17550 34783 17870 34784
rect 28620 34848 28940 34849
rect 28620 34784 28628 34848
rect 28692 34784 28708 34848
rect 28772 34784 28788 34848
rect 28852 34784 28868 34848
rect 28932 34784 28940 34848
rect 28620 34783 28940 34784
rect 12014 34304 12334 34305
rect 12014 34240 12022 34304
rect 12086 34240 12102 34304
rect 12166 34240 12182 34304
rect 12246 34240 12262 34304
rect 12326 34240 12334 34304
rect 12014 34239 12334 34240
rect 23085 34304 23405 34305
rect 23085 34240 23093 34304
rect 23157 34240 23173 34304
rect 23237 34240 23253 34304
rect 23317 34240 23333 34304
rect 23397 34240 23405 34304
rect 23085 34239 23405 34240
rect 6479 33760 6799 33761
rect 6479 33696 6487 33760
rect 6551 33696 6567 33760
rect 6631 33696 6647 33760
rect 6711 33696 6727 33760
rect 6791 33696 6799 33760
rect 6479 33695 6799 33696
rect 17550 33760 17870 33761
rect 17550 33696 17558 33760
rect 17622 33696 17638 33760
rect 17702 33696 17718 33760
rect 17782 33696 17798 33760
rect 17862 33696 17870 33760
rect 17550 33695 17870 33696
rect 28620 33760 28940 33761
rect 28620 33696 28628 33760
rect 28692 33696 28708 33760
rect 28772 33696 28788 33760
rect 28852 33696 28868 33760
rect 28932 33696 28940 33760
rect 28620 33695 28940 33696
rect 33593 33418 33659 33421
rect 34709 33418 35509 33448
rect 33593 33416 35509 33418
rect 33593 33360 33598 33416
rect 33654 33360 35509 33416
rect 33593 33358 35509 33360
rect 33593 33355 33659 33358
rect 34709 33328 35509 33358
rect 12014 33216 12334 33217
rect 12014 33152 12022 33216
rect 12086 33152 12102 33216
rect 12166 33152 12182 33216
rect 12246 33152 12262 33216
rect 12326 33152 12334 33216
rect 12014 33151 12334 33152
rect 23085 33216 23405 33217
rect 23085 33152 23093 33216
rect 23157 33152 23173 33216
rect 23237 33152 23253 33216
rect 23317 33152 23333 33216
rect 23397 33152 23405 33216
rect 23085 33151 23405 33152
rect 0 32738 800 32768
rect 1393 32738 1459 32741
rect 0 32736 1459 32738
rect 0 32680 1398 32736
rect 1454 32680 1459 32736
rect 0 32678 1459 32680
rect 0 32648 800 32678
rect 1393 32675 1459 32678
rect 6479 32672 6799 32673
rect 6479 32608 6487 32672
rect 6551 32608 6567 32672
rect 6631 32608 6647 32672
rect 6711 32608 6727 32672
rect 6791 32608 6799 32672
rect 6479 32607 6799 32608
rect 17550 32672 17870 32673
rect 17550 32608 17558 32672
rect 17622 32608 17638 32672
rect 17702 32608 17718 32672
rect 17782 32608 17798 32672
rect 17862 32608 17870 32672
rect 17550 32607 17870 32608
rect 28620 32672 28940 32673
rect 28620 32608 28628 32672
rect 28692 32608 28708 32672
rect 28772 32608 28788 32672
rect 28852 32608 28868 32672
rect 28932 32608 28940 32672
rect 28620 32607 28940 32608
rect 12014 32128 12334 32129
rect 12014 32064 12022 32128
rect 12086 32064 12102 32128
rect 12166 32064 12182 32128
rect 12246 32064 12262 32128
rect 12326 32064 12334 32128
rect 12014 32063 12334 32064
rect 23085 32128 23405 32129
rect 23085 32064 23093 32128
rect 23157 32064 23173 32128
rect 23237 32064 23253 32128
rect 23317 32064 23333 32128
rect 23397 32064 23405 32128
rect 23085 32063 23405 32064
rect 6479 31584 6799 31585
rect 6479 31520 6487 31584
rect 6551 31520 6567 31584
rect 6631 31520 6647 31584
rect 6711 31520 6727 31584
rect 6791 31520 6799 31584
rect 6479 31519 6799 31520
rect 17550 31584 17870 31585
rect 17550 31520 17558 31584
rect 17622 31520 17638 31584
rect 17702 31520 17718 31584
rect 17782 31520 17798 31584
rect 17862 31520 17870 31584
rect 17550 31519 17870 31520
rect 28620 31584 28940 31585
rect 28620 31520 28628 31584
rect 28692 31520 28708 31584
rect 28772 31520 28788 31584
rect 28852 31520 28868 31584
rect 28932 31520 28940 31584
rect 28620 31519 28940 31520
rect 12014 31040 12334 31041
rect 12014 30976 12022 31040
rect 12086 30976 12102 31040
rect 12166 30976 12182 31040
rect 12246 30976 12262 31040
rect 12326 30976 12334 31040
rect 12014 30975 12334 30976
rect 23085 31040 23405 31041
rect 23085 30976 23093 31040
rect 23157 30976 23173 31040
rect 23237 30976 23253 31040
rect 23317 30976 23333 31040
rect 23397 30976 23405 31040
rect 23085 30975 23405 30976
rect 6479 30496 6799 30497
rect 6479 30432 6487 30496
rect 6551 30432 6567 30496
rect 6631 30432 6647 30496
rect 6711 30432 6727 30496
rect 6791 30432 6799 30496
rect 6479 30431 6799 30432
rect 17550 30496 17870 30497
rect 17550 30432 17558 30496
rect 17622 30432 17638 30496
rect 17702 30432 17718 30496
rect 17782 30432 17798 30496
rect 17862 30432 17870 30496
rect 17550 30431 17870 30432
rect 28620 30496 28940 30497
rect 28620 30432 28628 30496
rect 28692 30432 28708 30496
rect 28772 30432 28788 30496
rect 28852 30432 28868 30496
rect 28932 30432 28940 30496
rect 28620 30431 28940 30432
rect 12014 29952 12334 29953
rect 12014 29888 12022 29952
rect 12086 29888 12102 29952
rect 12166 29888 12182 29952
rect 12246 29888 12262 29952
rect 12326 29888 12334 29952
rect 12014 29887 12334 29888
rect 23085 29952 23405 29953
rect 23085 29888 23093 29952
rect 23157 29888 23173 29952
rect 23237 29888 23253 29952
rect 23317 29888 23333 29952
rect 23397 29888 23405 29952
rect 23085 29887 23405 29888
rect 6479 29408 6799 29409
rect 6479 29344 6487 29408
rect 6551 29344 6567 29408
rect 6631 29344 6647 29408
rect 6711 29344 6727 29408
rect 6791 29344 6799 29408
rect 6479 29343 6799 29344
rect 17550 29408 17870 29409
rect 17550 29344 17558 29408
rect 17622 29344 17638 29408
rect 17702 29344 17718 29408
rect 17782 29344 17798 29408
rect 17862 29344 17870 29408
rect 17550 29343 17870 29344
rect 28620 29408 28940 29409
rect 28620 29344 28628 29408
rect 28692 29344 28708 29408
rect 28772 29344 28788 29408
rect 28852 29344 28868 29408
rect 28932 29344 28940 29408
rect 28620 29343 28940 29344
rect 33593 29338 33659 29341
rect 34709 29338 35509 29368
rect 33593 29336 35509 29338
rect 33593 29280 33598 29336
rect 33654 29280 35509 29336
rect 33593 29278 35509 29280
rect 33593 29275 33659 29278
rect 34709 29248 35509 29278
rect 12014 28864 12334 28865
rect 12014 28800 12022 28864
rect 12086 28800 12102 28864
rect 12166 28800 12182 28864
rect 12246 28800 12262 28864
rect 12326 28800 12334 28864
rect 12014 28799 12334 28800
rect 23085 28864 23405 28865
rect 23085 28800 23093 28864
rect 23157 28800 23173 28864
rect 23237 28800 23253 28864
rect 23317 28800 23333 28864
rect 23397 28800 23405 28864
rect 23085 28799 23405 28800
rect 0 28658 800 28688
rect 1761 28658 1827 28661
rect 0 28656 1827 28658
rect 0 28600 1766 28656
rect 1822 28600 1827 28656
rect 0 28598 1827 28600
rect 0 28568 800 28598
rect 1761 28595 1827 28598
rect 6479 28320 6799 28321
rect 6479 28256 6487 28320
rect 6551 28256 6567 28320
rect 6631 28256 6647 28320
rect 6711 28256 6727 28320
rect 6791 28256 6799 28320
rect 6479 28255 6799 28256
rect 17550 28320 17870 28321
rect 17550 28256 17558 28320
rect 17622 28256 17638 28320
rect 17702 28256 17718 28320
rect 17782 28256 17798 28320
rect 17862 28256 17870 28320
rect 17550 28255 17870 28256
rect 28620 28320 28940 28321
rect 28620 28256 28628 28320
rect 28692 28256 28708 28320
rect 28772 28256 28788 28320
rect 28852 28256 28868 28320
rect 28932 28256 28940 28320
rect 28620 28255 28940 28256
rect 12014 27776 12334 27777
rect 12014 27712 12022 27776
rect 12086 27712 12102 27776
rect 12166 27712 12182 27776
rect 12246 27712 12262 27776
rect 12326 27712 12334 27776
rect 12014 27711 12334 27712
rect 23085 27776 23405 27777
rect 23085 27712 23093 27776
rect 23157 27712 23173 27776
rect 23237 27712 23253 27776
rect 23317 27712 23333 27776
rect 23397 27712 23405 27776
rect 23085 27711 23405 27712
rect 6479 27232 6799 27233
rect 6479 27168 6487 27232
rect 6551 27168 6567 27232
rect 6631 27168 6647 27232
rect 6711 27168 6727 27232
rect 6791 27168 6799 27232
rect 6479 27167 6799 27168
rect 17550 27232 17870 27233
rect 17550 27168 17558 27232
rect 17622 27168 17638 27232
rect 17702 27168 17718 27232
rect 17782 27168 17798 27232
rect 17862 27168 17870 27232
rect 17550 27167 17870 27168
rect 28620 27232 28940 27233
rect 28620 27168 28628 27232
rect 28692 27168 28708 27232
rect 28772 27168 28788 27232
rect 28852 27168 28868 27232
rect 28932 27168 28940 27232
rect 28620 27167 28940 27168
rect 12014 26688 12334 26689
rect 12014 26624 12022 26688
rect 12086 26624 12102 26688
rect 12166 26624 12182 26688
rect 12246 26624 12262 26688
rect 12326 26624 12334 26688
rect 12014 26623 12334 26624
rect 23085 26688 23405 26689
rect 23085 26624 23093 26688
rect 23157 26624 23173 26688
rect 23237 26624 23253 26688
rect 23317 26624 23333 26688
rect 23397 26624 23405 26688
rect 23085 26623 23405 26624
rect 6479 26144 6799 26145
rect 6479 26080 6487 26144
rect 6551 26080 6567 26144
rect 6631 26080 6647 26144
rect 6711 26080 6727 26144
rect 6791 26080 6799 26144
rect 6479 26079 6799 26080
rect 17550 26144 17870 26145
rect 17550 26080 17558 26144
rect 17622 26080 17638 26144
rect 17702 26080 17718 26144
rect 17782 26080 17798 26144
rect 17862 26080 17870 26144
rect 17550 26079 17870 26080
rect 28620 26144 28940 26145
rect 28620 26080 28628 26144
rect 28692 26080 28708 26144
rect 28772 26080 28788 26144
rect 28852 26080 28868 26144
rect 28932 26080 28940 26144
rect 28620 26079 28940 26080
rect 12014 25600 12334 25601
rect 12014 25536 12022 25600
rect 12086 25536 12102 25600
rect 12166 25536 12182 25600
rect 12246 25536 12262 25600
rect 12326 25536 12334 25600
rect 12014 25535 12334 25536
rect 23085 25600 23405 25601
rect 23085 25536 23093 25600
rect 23157 25536 23173 25600
rect 23237 25536 23253 25600
rect 23317 25536 23333 25600
rect 23397 25536 23405 25600
rect 23085 25535 23405 25536
rect 11145 25394 11211 25397
rect 12801 25394 12867 25397
rect 11145 25392 12867 25394
rect 11145 25336 11150 25392
rect 11206 25336 12806 25392
rect 12862 25336 12867 25392
rect 11145 25334 12867 25336
rect 11145 25331 11211 25334
rect 12801 25331 12867 25334
rect 33501 25258 33567 25261
rect 34709 25258 35509 25288
rect 33501 25256 35509 25258
rect 33501 25200 33506 25256
rect 33562 25200 35509 25256
rect 33501 25198 35509 25200
rect 33501 25195 33567 25198
rect 34709 25168 35509 25198
rect 6479 25056 6799 25057
rect 6479 24992 6487 25056
rect 6551 24992 6567 25056
rect 6631 24992 6647 25056
rect 6711 24992 6727 25056
rect 6791 24992 6799 25056
rect 6479 24991 6799 24992
rect 17550 25056 17870 25057
rect 17550 24992 17558 25056
rect 17622 24992 17638 25056
rect 17702 24992 17718 25056
rect 17782 24992 17798 25056
rect 17862 24992 17870 25056
rect 17550 24991 17870 24992
rect 28620 25056 28940 25057
rect 28620 24992 28628 25056
rect 28692 24992 28708 25056
rect 28772 24992 28788 25056
rect 28852 24992 28868 25056
rect 28932 24992 28940 25056
rect 28620 24991 28940 24992
rect 0 24578 800 24608
rect 1393 24578 1459 24581
rect 0 24576 1459 24578
rect 0 24520 1398 24576
rect 1454 24520 1459 24576
rect 0 24518 1459 24520
rect 0 24488 800 24518
rect 1393 24515 1459 24518
rect 12014 24512 12334 24513
rect 12014 24448 12022 24512
rect 12086 24448 12102 24512
rect 12166 24448 12182 24512
rect 12246 24448 12262 24512
rect 12326 24448 12334 24512
rect 12014 24447 12334 24448
rect 23085 24512 23405 24513
rect 23085 24448 23093 24512
rect 23157 24448 23173 24512
rect 23237 24448 23253 24512
rect 23317 24448 23333 24512
rect 23397 24448 23405 24512
rect 23085 24447 23405 24448
rect 6479 23968 6799 23969
rect 6479 23904 6487 23968
rect 6551 23904 6567 23968
rect 6631 23904 6647 23968
rect 6711 23904 6727 23968
rect 6791 23904 6799 23968
rect 6479 23903 6799 23904
rect 17550 23968 17870 23969
rect 17550 23904 17558 23968
rect 17622 23904 17638 23968
rect 17702 23904 17718 23968
rect 17782 23904 17798 23968
rect 17862 23904 17870 23968
rect 17550 23903 17870 23904
rect 28620 23968 28940 23969
rect 28620 23904 28628 23968
rect 28692 23904 28708 23968
rect 28772 23904 28788 23968
rect 28852 23904 28868 23968
rect 28932 23904 28940 23968
rect 28620 23903 28940 23904
rect 12014 23424 12334 23425
rect 12014 23360 12022 23424
rect 12086 23360 12102 23424
rect 12166 23360 12182 23424
rect 12246 23360 12262 23424
rect 12326 23360 12334 23424
rect 12014 23359 12334 23360
rect 23085 23424 23405 23425
rect 23085 23360 23093 23424
rect 23157 23360 23173 23424
rect 23237 23360 23253 23424
rect 23317 23360 23333 23424
rect 23397 23360 23405 23424
rect 23085 23359 23405 23360
rect 6479 22880 6799 22881
rect 6479 22816 6487 22880
rect 6551 22816 6567 22880
rect 6631 22816 6647 22880
rect 6711 22816 6727 22880
rect 6791 22816 6799 22880
rect 6479 22815 6799 22816
rect 17550 22880 17870 22881
rect 17550 22816 17558 22880
rect 17622 22816 17638 22880
rect 17702 22816 17718 22880
rect 17782 22816 17798 22880
rect 17862 22816 17870 22880
rect 17550 22815 17870 22816
rect 28620 22880 28940 22881
rect 28620 22816 28628 22880
rect 28692 22816 28708 22880
rect 28772 22816 28788 22880
rect 28852 22816 28868 22880
rect 28932 22816 28940 22880
rect 28620 22815 28940 22816
rect 12014 22336 12334 22337
rect 12014 22272 12022 22336
rect 12086 22272 12102 22336
rect 12166 22272 12182 22336
rect 12246 22272 12262 22336
rect 12326 22272 12334 22336
rect 12014 22271 12334 22272
rect 23085 22336 23405 22337
rect 23085 22272 23093 22336
rect 23157 22272 23173 22336
rect 23237 22272 23253 22336
rect 23317 22272 23333 22336
rect 23397 22272 23405 22336
rect 23085 22271 23405 22272
rect 12157 21994 12223 21997
rect 16573 21994 16639 21997
rect 12157 21992 16639 21994
rect 12157 21936 12162 21992
rect 12218 21936 16578 21992
rect 16634 21936 16639 21992
rect 12157 21934 16639 21936
rect 12157 21931 12223 21934
rect 16573 21931 16639 21934
rect 6479 21792 6799 21793
rect 6479 21728 6487 21792
rect 6551 21728 6567 21792
rect 6631 21728 6647 21792
rect 6711 21728 6727 21792
rect 6791 21728 6799 21792
rect 6479 21727 6799 21728
rect 17550 21792 17870 21793
rect 17550 21728 17558 21792
rect 17622 21728 17638 21792
rect 17702 21728 17718 21792
rect 17782 21728 17798 21792
rect 17862 21728 17870 21792
rect 17550 21727 17870 21728
rect 28620 21792 28940 21793
rect 28620 21728 28628 21792
rect 28692 21728 28708 21792
rect 28772 21728 28788 21792
rect 28852 21728 28868 21792
rect 28932 21728 28940 21792
rect 28620 21727 28940 21728
rect 12014 21248 12334 21249
rect 12014 21184 12022 21248
rect 12086 21184 12102 21248
rect 12166 21184 12182 21248
rect 12246 21184 12262 21248
rect 12326 21184 12334 21248
rect 12014 21183 12334 21184
rect 23085 21248 23405 21249
rect 23085 21184 23093 21248
rect 23157 21184 23173 21248
rect 23237 21184 23253 21248
rect 23317 21184 23333 21248
rect 23397 21184 23405 21248
rect 23085 21183 23405 21184
rect 33593 21178 33659 21181
rect 34709 21178 35509 21208
rect 33593 21176 35509 21178
rect 33593 21120 33598 21176
rect 33654 21120 35509 21176
rect 33593 21118 35509 21120
rect 33593 21115 33659 21118
rect 34709 21088 35509 21118
rect 6479 20704 6799 20705
rect 6479 20640 6487 20704
rect 6551 20640 6567 20704
rect 6631 20640 6647 20704
rect 6711 20640 6727 20704
rect 6791 20640 6799 20704
rect 6479 20639 6799 20640
rect 17550 20704 17870 20705
rect 17550 20640 17558 20704
rect 17622 20640 17638 20704
rect 17702 20640 17718 20704
rect 17782 20640 17798 20704
rect 17862 20640 17870 20704
rect 17550 20639 17870 20640
rect 28620 20704 28940 20705
rect 28620 20640 28628 20704
rect 28692 20640 28708 20704
rect 28772 20640 28788 20704
rect 28852 20640 28868 20704
rect 28932 20640 28940 20704
rect 28620 20639 28940 20640
rect 0 20498 800 20528
rect 1761 20498 1827 20501
rect 0 20496 1827 20498
rect 0 20440 1766 20496
rect 1822 20440 1827 20496
rect 0 20438 1827 20440
rect 0 20408 800 20438
rect 1761 20435 1827 20438
rect 12014 20160 12334 20161
rect 12014 20096 12022 20160
rect 12086 20096 12102 20160
rect 12166 20096 12182 20160
rect 12246 20096 12262 20160
rect 12326 20096 12334 20160
rect 12014 20095 12334 20096
rect 23085 20160 23405 20161
rect 23085 20096 23093 20160
rect 23157 20096 23173 20160
rect 23237 20096 23253 20160
rect 23317 20096 23333 20160
rect 23397 20096 23405 20160
rect 23085 20095 23405 20096
rect 6479 19616 6799 19617
rect 6479 19552 6487 19616
rect 6551 19552 6567 19616
rect 6631 19552 6647 19616
rect 6711 19552 6727 19616
rect 6791 19552 6799 19616
rect 6479 19551 6799 19552
rect 17550 19616 17870 19617
rect 17550 19552 17558 19616
rect 17622 19552 17638 19616
rect 17702 19552 17718 19616
rect 17782 19552 17798 19616
rect 17862 19552 17870 19616
rect 17550 19551 17870 19552
rect 28620 19616 28940 19617
rect 28620 19552 28628 19616
rect 28692 19552 28708 19616
rect 28772 19552 28788 19616
rect 28852 19552 28868 19616
rect 28932 19552 28940 19616
rect 28620 19551 28940 19552
rect 20621 19410 20687 19413
rect 22461 19410 22527 19413
rect 20621 19408 22527 19410
rect 20621 19352 20626 19408
rect 20682 19352 22466 19408
rect 22522 19352 22527 19408
rect 20621 19350 22527 19352
rect 20621 19347 20687 19350
rect 22461 19347 22527 19350
rect 13353 19274 13419 19277
rect 14641 19274 14707 19277
rect 13353 19272 14707 19274
rect 13353 19216 13358 19272
rect 13414 19216 14646 19272
rect 14702 19216 14707 19272
rect 13353 19214 14707 19216
rect 13353 19211 13419 19214
rect 14641 19211 14707 19214
rect 15009 19274 15075 19277
rect 17309 19274 17375 19277
rect 15009 19272 17375 19274
rect 15009 19216 15014 19272
rect 15070 19216 17314 19272
rect 17370 19216 17375 19272
rect 15009 19214 17375 19216
rect 15009 19211 15075 19214
rect 17309 19211 17375 19214
rect 12014 19072 12334 19073
rect 12014 19008 12022 19072
rect 12086 19008 12102 19072
rect 12166 19008 12182 19072
rect 12246 19008 12262 19072
rect 12326 19008 12334 19072
rect 12014 19007 12334 19008
rect 23085 19072 23405 19073
rect 23085 19008 23093 19072
rect 23157 19008 23173 19072
rect 23237 19008 23253 19072
rect 23317 19008 23333 19072
rect 23397 19008 23405 19072
rect 23085 19007 23405 19008
rect 19885 18866 19951 18869
rect 25589 18866 25655 18869
rect 19885 18864 25655 18866
rect 19885 18808 19890 18864
rect 19946 18808 25594 18864
rect 25650 18808 25655 18864
rect 19885 18806 25655 18808
rect 19885 18803 19951 18806
rect 25589 18803 25655 18806
rect 12249 18594 12315 18597
rect 16665 18594 16731 18597
rect 12249 18592 16731 18594
rect 12249 18536 12254 18592
rect 12310 18536 16670 18592
rect 16726 18536 16731 18592
rect 12249 18534 16731 18536
rect 12249 18531 12315 18534
rect 16665 18531 16731 18534
rect 6479 18528 6799 18529
rect 6479 18464 6487 18528
rect 6551 18464 6567 18528
rect 6631 18464 6647 18528
rect 6711 18464 6727 18528
rect 6791 18464 6799 18528
rect 6479 18463 6799 18464
rect 17550 18528 17870 18529
rect 17550 18464 17558 18528
rect 17622 18464 17638 18528
rect 17702 18464 17718 18528
rect 17782 18464 17798 18528
rect 17862 18464 17870 18528
rect 17550 18463 17870 18464
rect 28620 18528 28940 18529
rect 28620 18464 28628 18528
rect 28692 18464 28708 18528
rect 28772 18464 28788 18528
rect 28852 18464 28868 18528
rect 28932 18464 28940 18528
rect 28620 18463 28940 18464
rect 12014 17984 12334 17985
rect 12014 17920 12022 17984
rect 12086 17920 12102 17984
rect 12166 17920 12182 17984
rect 12246 17920 12262 17984
rect 12326 17920 12334 17984
rect 12014 17919 12334 17920
rect 23085 17984 23405 17985
rect 23085 17920 23093 17984
rect 23157 17920 23173 17984
rect 23237 17920 23253 17984
rect 23317 17920 23333 17984
rect 23397 17920 23405 17984
rect 23085 17919 23405 17920
rect 6479 17440 6799 17441
rect 6479 17376 6487 17440
rect 6551 17376 6567 17440
rect 6631 17376 6647 17440
rect 6711 17376 6727 17440
rect 6791 17376 6799 17440
rect 6479 17375 6799 17376
rect 17550 17440 17870 17441
rect 17550 17376 17558 17440
rect 17622 17376 17638 17440
rect 17702 17376 17718 17440
rect 17782 17376 17798 17440
rect 17862 17376 17870 17440
rect 17550 17375 17870 17376
rect 28620 17440 28940 17441
rect 28620 17376 28628 17440
rect 28692 17376 28708 17440
rect 28772 17376 28788 17440
rect 28852 17376 28868 17440
rect 28932 17376 28940 17440
rect 28620 17375 28940 17376
rect 33593 17098 33659 17101
rect 34709 17098 35509 17128
rect 33593 17096 35509 17098
rect 33593 17040 33598 17096
rect 33654 17040 35509 17096
rect 33593 17038 35509 17040
rect 33593 17035 33659 17038
rect 34709 17008 35509 17038
rect 12014 16896 12334 16897
rect 12014 16832 12022 16896
rect 12086 16832 12102 16896
rect 12166 16832 12182 16896
rect 12246 16832 12262 16896
rect 12326 16832 12334 16896
rect 12014 16831 12334 16832
rect 23085 16896 23405 16897
rect 23085 16832 23093 16896
rect 23157 16832 23173 16896
rect 23237 16832 23253 16896
rect 23317 16832 23333 16896
rect 23397 16832 23405 16896
rect 23085 16831 23405 16832
rect 0 16418 800 16448
rect 4061 16418 4127 16421
rect 0 16416 4127 16418
rect 0 16360 4066 16416
rect 4122 16360 4127 16416
rect 0 16358 4127 16360
rect 0 16328 800 16358
rect 4061 16355 4127 16358
rect 6479 16352 6799 16353
rect 6479 16288 6487 16352
rect 6551 16288 6567 16352
rect 6631 16288 6647 16352
rect 6711 16288 6727 16352
rect 6791 16288 6799 16352
rect 6479 16287 6799 16288
rect 17550 16352 17870 16353
rect 17550 16288 17558 16352
rect 17622 16288 17638 16352
rect 17702 16288 17718 16352
rect 17782 16288 17798 16352
rect 17862 16288 17870 16352
rect 17550 16287 17870 16288
rect 28620 16352 28940 16353
rect 28620 16288 28628 16352
rect 28692 16288 28708 16352
rect 28772 16288 28788 16352
rect 28852 16288 28868 16352
rect 28932 16288 28940 16352
rect 28620 16287 28940 16288
rect 12014 15808 12334 15809
rect 12014 15744 12022 15808
rect 12086 15744 12102 15808
rect 12166 15744 12182 15808
rect 12246 15744 12262 15808
rect 12326 15744 12334 15808
rect 12014 15743 12334 15744
rect 23085 15808 23405 15809
rect 23085 15744 23093 15808
rect 23157 15744 23173 15808
rect 23237 15744 23253 15808
rect 23317 15744 23333 15808
rect 23397 15744 23405 15808
rect 23085 15743 23405 15744
rect 6479 15264 6799 15265
rect 6479 15200 6487 15264
rect 6551 15200 6567 15264
rect 6631 15200 6647 15264
rect 6711 15200 6727 15264
rect 6791 15200 6799 15264
rect 6479 15199 6799 15200
rect 17550 15264 17870 15265
rect 17550 15200 17558 15264
rect 17622 15200 17638 15264
rect 17702 15200 17718 15264
rect 17782 15200 17798 15264
rect 17862 15200 17870 15264
rect 17550 15199 17870 15200
rect 28620 15264 28940 15265
rect 28620 15200 28628 15264
rect 28692 15200 28708 15264
rect 28772 15200 28788 15264
rect 28852 15200 28868 15264
rect 28932 15200 28940 15264
rect 28620 15199 28940 15200
rect 12014 14720 12334 14721
rect 12014 14656 12022 14720
rect 12086 14656 12102 14720
rect 12166 14656 12182 14720
rect 12246 14656 12262 14720
rect 12326 14656 12334 14720
rect 12014 14655 12334 14656
rect 23085 14720 23405 14721
rect 23085 14656 23093 14720
rect 23157 14656 23173 14720
rect 23237 14656 23253 14720
rect 23317 14656 23333 14720
rect 23397 14656 23405 14720
rect 23085 14655 23405 14656
rect 6479 14176 6799 14177
rect 6479 14112 6487 14176
rect 6551 14112 6567 14176
rect 6631 14112 6647 14176
rect 6711 14112 6727 14176
rect 6791 14112 6799 14176
rect 6479 14111 6799 14112
rect 17550 14176 17870 14177
rect 17550 14112 17558 14176
rect 17622 14112 17638 14176
rect 17702 14112 17718 14176
rect 17782 14112 17798 14176
rect 17862 14112 17870 14176
rect 17550 14111 17870 14112
rect 28620 14176 28940 14177
rect 28620 14112 28628 14176
rect 28692 14112 28708 14176
rect 28772 14112 28788 14176
rect 28852 14112 28868 14176
rect 28932 14112 28940 14176
rect 28620 14111 28940 14112
rect 12014 13632 12334 13633
rect 12014 13568 12022 13632
rect 12086 13568 12102 13632
rect 12166 13568 12182 13632
rect 12246 13568 12262 13632
rect 12326 13568 12334 13632
rect 12014 13567 12334 13568
rect 23085 13632 23405 13633
rect 23085 13568 23093 13632
rect 23157 13568 23173 13632
rect 23237 13568 23253 13632
rect 23317 13568 23333 13632
rect 23397 13568 23405 13632
rect 23085 13567 23405 13568
rect 6479 13088 6799 13089
rect 6479 13024 6487 13088
rect 6551 13024 6567 13088
rect 6631 13024 6647 13088
rect 6711 13024 6727 13088
rect 6791 13024 6799 13088
rect 6479 13023 6799 13024
rect 17550 13088 17870 13089
rect 17550 13024 17558 13088
rect 17622 13024 17638 13088
rect 17702 13024 17718 13088
rect 17782 13024 17798 13088
rect 17862 13024 17870 13088
rect 17550 13023 17870 13024
rect 28620 13088 28940 13089
rect 28620 13024 28628 13088
rect 28692 13024 28708 13088
rect 28772 13024 28788 13088
rect 28852 13024 28868 13088
rect 28932 13024 28940 13088
rect 28620 13023 28940 13024
rect 33593 13018 33659 13021
rect 34709 13018 35509 13048
rect 33593 13016 35509 13018
rect 33593 12960 33598 13016
rect 33654 12960 35509 13016
rect 33593 12958 35509 12960
rect 33593 12955 33659 12958
rect 34709 12928 35509 12958
rect 12014 12544 12334 12545
rect 12014 12480 12022 12544
rect 12086 12480 12102 12544
rect 12166 12480 12182 12544
rect 12246 12480 12262 12544
rect 12326 12480 12334 12544
rect 12014 12479 12334 12480
rect 23085 12544 23405 12545
rect 23085 12480 23093 12544
rect 23157 12480 23173 12544
rect 23237 12480 23253 12544
rect 23317 12480 23333 12544
rect 23397 12480 23405 12544
rect 23085 12479 23405 12480
rect 0 12338 800 12368
rect 1761 12338 1827 12341
rect 0 12336 1827 12338
rect 0 12280 1766 12336
rect 1822 12280 1827 12336
rect 0 12278 1827 12280
rect 0 12248 800 12278
rect 1761 12275 1827 12278
rect 6479 12000 6799 12001
rect 6479 11936 6487 12000
rect 6551 11936 6567 12000
rect 6631 11936 6647 12000
rect 6711 11936 6727 12000
rect 6791 11936 6799 12000
rect 6479 11935 6799 11936
rect 17550 12000 17870 12001
rect 17550 11936 17558 12000
rect 17622 11936 17638 12000
rect 17702 11936 17718 12000
rect 17782 11936 17798 12000
rect 17862 11936 17870 12000
rect 17550 11935 17870 11936
rect 28620 12000 28940 12001
rect 28620 11936 28628 12000
rect 28692 11936 28708 12000
rect 28772 11936 28788 12000
rect 28852 11936 28868 12000
rect 28932 11936 28940 12000
rect 28620 11935 28940 11936
rect 12014 11456 12334 11457
rect 12014 11392 12022 11456
rect 12086 11392 12102 11456
rect 12166 11392 12182 11456
rect 12246 11392 12262 11456
rect 12326 11392 12334 11456
rect 12014 11391 12334 11392
rect 23085 11456 23405 11457
rect 23085 11392 23093 11456
rect 23157 11392 23173 11456
rect 23237 11392 23253 11456
rect 23317 11392 23333 11456
rect 23397 11392 23405 11456
rect 23085 11391 23405 11392
rect 6479 10912 6799 10913
rect 6479 10848 6487 10912
rect 6551 10848 6567 10912
rect 6631 10848 6647 10912
rect 6711 10848 6727 10912
rect 6791 10848 6799 10912
rect 6479 10847 6799 10848
rect 17550 10912 17870 10913
rect 17550 10848 17558 10912
rect 17622 10848 17638 10912
rect 17702 10848 17718 10912
rect 17782 10848 17798 10912
rect 17862 10848 17870 10912
rect 17550 10847 17870 10848
rect 28620 10912 28940 10913
rect 28620 10848 28628 10912
rect 28692 10848 28708 10912
rect 28772 10848 28788 10912
rect 28852 10848 28868 10912
rect 28932 10848 28940 10912
rect 28620 10847 28940 10848
rect 12014 10368 12334 10369
rect 12014 10304 12022 10368
rect 12086 10304 12102 10368
rect 12166 10304 12182 10368
rect 12246 10304 12262 10368
rect 12326 10304 12334 10368
rect 12014 10303 12334 10304
rect 23085 10368 23405 10369
rect 23085 10304 23093 10368
rect 23157 10304 23173 10368
rect 23237 10304 23253 10368
rect 23317 10304 23333 10368
rect 23397 10304 23405 10368
rect 23085 10303 23405 10304
rect 6479 9824 6799 9825
rect 6479 9760 6487 9824
rect 6551 9760 6567 9824
rect 6631 9760 6647 9824
rect 6711 9760 6727 9824
rect 6791 9760 6799 9824
rect 6479 9759 6799 9760
rect 17550 9824 17870 9825
rect 17550 9760 17558 9824
rect 17622 9760 17638 9824
rect 17702 9760 17718 9824
rect 17782 9760 17798 9824
rect 17862 9760 17870 9824
rect 17550 9759 17870 9760
rect 28620 9824 28940 9825
rect 28620 9760 28628 9824
rect 28692 9760 28708 9824
rect 28772 9760 28788 9824
rect 28852 9760 28868 9824
rect 28932 9760 28940 9824
rect 28620 9759 28940 9760
rect 12014 9280 12334 9281
rect 12014 9216 12022 9280
rect 12086 9216 12102 9280
rect 12166 9216 12182 9280
rect 12246 9216 12262 9280
rect 12326 9216 12334 9280
rect 12014 9215 12334 9216
rect 23085 9280 23405 9281
rect 23085 9216 23093 9280
rect 23157 9216 23173 9280
rect 23237 9216 23253 9280
rect 23317 9216 23333 9280
rect 23397 9216 23405 9280
rect 23085 9215 23405 9216
rect 30465 8938 30531 8941
rect 34709 8938 35509 8968
rect 30465 8936 35509 8938
rect 30465 8880 30470 8936
rect 30526 8880 35509 8936
rect 30465 8878 35509 8880
rect 30465 8875 30531 8878
rect 34709 8848 35509 8878
rect 6479 8736 6799 8737
rect 6479 8672 6487 8736
rect 6551 8672 6567 8736
rect 6631 8672 6647 8736
rect 6711 8672 6727 8736
rect 6791 8672 6799 8736
rect 6479 8671 6799 8672
rect 17550 8736 17870 8737
rect 17550 8672 17558 8736
rect 17622 8672 17638 8736
rect 17702 8672 17718 8736
rect 17782 8672 17798 8736
rect 17862 8672 17870 8736
rect 17550 8671 17870 8672
rect 28620 8736 28940 8737
rect 28620 8672 28628 8736
rect 28692 8672 28708 8736
rect 28772 8672 28788 8736
rect 28852 8672 28868 8736
rect 28932 8672 28940 8736
rect 28620 8671 28940 8672
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 12014 8192 12334 8193
rect 12014 8128 12022 8192
rect 12086 8128 12102 8192
rect 12166 8128 12182 8192
rect 12246 8128 12262 8192
rect 12326 8128 12334 8192
rect 12014 8127 12334 8128
rect 23085 8192 23405 8193
rect 23085 8128 23093 8192
rect 23157 8128 23173 8192
rect 23237 8128 23253 8192
rect 23317 8128 23333 8192
rect 23397 8128 23405 8192
rect 23085 8127 23405 8128
rect 6479 7648 6799 7649
rect 6479 7584 6487 7648
rect 6551 7584 6567 7648
rect 6631 7584 6647 7648
rect 6711 7584 6727 7648
rect 6791 7584 6799 7648
rect 6479 7583 6799 7584
rect 17550 7648 17870 7649
rect 17550 7584 17558 7648
rect 17622 7584 17638 7648
rect 17702 7584 17718 7648
rect 17782 7584 17798 7648
rect 17862 7584 17870 7648
rect 17550 7583 17870 7584
rect 28620 7648 28940 7649
rect 28620 7584 28628 7648
rect 28692 7584 28708 7648
rect 28772 7584 28788 7648
rect 28852 7584 28868 7648
rect 28932 7584 28940 7648
rect 28620 7583 28940 7584
rect 12014 7104 12334 7105
rect 12014 7040 12022 7104
rect 12086 7040 12102 7104
rect 12166 7040 12182 7104
rect 12246 7040 12262 7104
rect 12326 7040 12334 7104
rect 12014 7039 12334 7040
rect 23085 7104 23405 7105
rect 23085 7040 23093 7104
rect 23157 7040 23173 7104
rect 23237 7040 23253 7104
rect 23317 7040 23333 7104
rect 23397 7040 23405 7104
rect 23085 7039 23405 7040
rect 6479 6560 6799 6561
rect 6479 6496 6487 6560
rect 6551 6496 6567 6560
rect 6631 6496 6647 6560
rect 6711 6496 6727 6560
rect 6791 6496 6799 6560
rect 6479 6495 6799 6496
rect 17550 6560 17870 6561
rect 17550 6496 17558 6560
rect 17622 6496 17638 6560
rect 17702 6496 17718 6560
rect 17782 6496 17798 6560
rect 17862 6496 17870 6560
rect 17550 6495 17870 6496
rect 28620 6560 28940 6561
rect 28620 6496 28628 6560
rect 28692 6496 28708 6560
rect 28772 6496 28788 6560
rect 28852 6496 28868 6560
rect 28932 6496 28940 6560
rect 28620 6495 28940 6496
rect 12014 6016 12334 6017
rect 12014 5952 12022 6016
rect 12086 5952 12102 6016
rect 12166 5952 12182 6016
rect 12246 5952 12262 6016
rect 12326 5952 12334 6016
rect 12014 5951 12334 5952
rect 23085 6016 23405 6017
rect 23085 5952 23093 6016
rect 23157 5952 23173 6016
rect 23237 5952 23253 6016
rect 23317 5952 23333 6016
rect 23397 5952 23405 6016
rect 23085 5951 23405 5952
rect 6479 5472 6799 5473
rect 6479 5408 6487 5472
rect 6551 5408 6567 5472
rect 6631 5408 6647 5472
rect 6711 5408 6727 5472
rect 6791 5408 6799 5472
rect 6479 5407 6799 5408
rect 17550 5472 17870 5473
rect 17550 5408 17558 5472
rect 17622 5408 17638 5472
rect 17702 5408 17718 5472
rect 17782 5408 17798 5472
rect 17862 5408 17870 5472
rect 17550 5407 17870 5408
rect 28620 5472 28940 5473
rect 28620 5408 28628 5472
rect 28692 5408 28708 5472
rect 28772 5408 28788 5472
rect 28852 5408 28868 5472
rect 28932 5408 28940 5472
rect 28620 5407 28940 5408
rect 12014 4928 12334 4929
rect 12014 4864 12022 4928
rect 12086 4864 12102 4928
rect 12166 4864 12182 4928
rect 12246 4864 12262 4928
rect 12326 4864 12334 4928
rect 12014 4863 12334 4864
rect 23085 4928 23405 4929
rect 23085 4864 23093 4928
rect 23157 4864 23173 4928
rect 23237 4864 23253 4928
rect 23317 4864 23333 4928
rect 23397 4864 23405 4928
rect 23085 4863 23405 4864
rect 33593 4858 33659 4861
rect 34709 4858 35509 4888
rect 33593 4856 35509 4858
rect 33593 4800 33598 4856
rect 33654 4800 35509 4856
rect 33593 4798 35509 4800
rect 33593 4795 33659 4798
rect 34709 4768 35509 4798
rect 6479 4384 6799 4385
rect 6479 4320 6487 4384
rect 6551 4320 6567 4384
rect 6631 4320 6647 4384
rect 6711 4320 6727 4384
rect 6791 4320 6799 4384
rect 6479 4319 6799 4320
rect 17550 4384 17870 4385
rect 17550 4320 17558 4384
rect 17622 4320 17638 4384
rect 17702 4320 17718 4384
rect 17782 4320 17798 4384
rect 17862 4320 17870 4384
rect 17550 4319 17870 4320
rect 28620 4384 28940 4385
rect 28620 4320 28628 4384
rect 28692 4320 28708 4384
rect 28772 4320 28788 4384
rect 28852 4320 28868 4384
rect 28932 4320 28940 4384
rect 28620 4319 28940 4320
rect 0 4178 800 4208
rect 1853 4178 1919 4181
rect 0 4176 1919 4178
rect 0 4120 1858 4176
rect 1914 4120 1919 4176
rect 0 4118 1919 4120
rect 0 4088 800 4118
rect 1853 4115 1919 4118
rect 12014 3840 12334 3841
rect 12014 3776 12022 3840
rect 12086 3776 12102 3840
rect 12166 3776 12182 3840
rect 12246 3776 12262 3840
rect 12326 3776 12334 3840
rect 12014 3775 12334 3776
rect 23085 3840 23405 3841
rect 23085 3776 23093 3840
rect 23157 3776 23173 3840
rect 23237 3776 23253 3840
rect 23317 3776 23333 3840
rect 23397 3776 23405 3840
rect 23085 3775 23405 3776
rect 6479 3296 6799 3297
rect 6479 3232 6487 3296
rect 6551 3232 6567 3296
rect 6631 3232 6647 3296
rect 6711 3232 6727 3296
rect 6791 3232 6799 3296
rect 6479 3231 6799 3232
rect 17550 3296 17870 3297
rect 17550 3232 17558 3296
rect 17622 3232 17638 3296
rect 17702 3232 17718 3296
rect 17782 3232 17798 3296
rect 17862 3232 17870 3296
rect 17550 3231 17870 3232
rect 28620 3296 28940 3297
rect 28620 3232 28628 3296
rect 28692 3232 28708 3296
rect 28772 3232 28788 3296
rect 28852 3232 28868 3296
rect 28932 3232 28940 3296
rect 28620 3231 28940 3232
rect 12014 2752 12334 2753
rect 12014 2688 12022 2752
rect 12086 2688 12102 2752
rect 12166 2688 12182 2752
rect 12246 2688 12262 2752
rect 12326 2688 12334 2752
rect 12014 2687 12334 2688
rect 23085 2752 23405 2753
rect 23085 2688 23093 2752
rect 23157 2688 23173 2752
rect 23237 2688 23253 2752
rect 23317 2688 23333 2752
rect 23397 2688 23405 2752
rect 23085 2687 23405 2688
rect 6479 2208 6799 2209
rect 6479 2144 6487 2208
rect 6551 2144 6567 2208
rect 6631 2144 6647 2208
rect 6711 2144 6727 2208
rect 6791 2144 6799 2208
rect 6479 2143 6799 2144
rect 17550 2208 17870 2209
rect 17550 2144 17558 2208
rect 17622 2144 17638 2208
rect 17702 2144 17718 2208
rect 17782 2144 17798 2208
rect 17862 2144 17870 2208
rect 17550 2143 17870 2144
rect 28620 2208 28940 2209
rect 28620 2144 28628 2208
rect 28692 2144 28708 2208
rect 28772 2144 28788 2208
rect 28852 2144 28868 2208
rect 28932 2144 28940 2208
rect 28620 2143 28940 2144
rect 31937 778 32003 781
rect 34709 778 35509 808
rect 31937 776 35509 778
rect 31937 720 31942 776
rect 31998 720 35509 776
rect 31937 718 35509 720
rect 31937 715 32003 718
rect 34709 688 35509 718
<< via3 >>
rect 12022 35388 12086 35392
rect 12022 35332 12026 35388
rect 12026 35332 12082 35388
rect 12082 35332 12086 35388
rect 12022 35328 12086 35332
rect 12102 35388 12166 35392
rect 12102 35332 12106 35388
rect 12106 35332 12162 35388
rect 12162 35332 12166 35388
rect 12102 35328 12166 35332
rect 12182 35388 12246 35392
rect 12182 35332 12186 35388
rect 12186 35332 12242 35388
rect 12242 35332 12246 35388
rect 12182 35328 12246 35332
rect 12262 35388 12326 35392
rect 12262 35332 12266 35388
rect 12266 35332 12322 35388
rect 12322 35332 12326 35388
rect 12262 35328 12326 35332
rect 23093 35388 23157 35392
rect 23093 35332 23097 35388
rect 23097 35332 23153 35388
rect 23153 35332 23157 35388
rect 23093 35328 23157 35332
rect 23173 35388 23237 35392
rect 23173 35332 23177 35388
rect 23177 35332 23233 35388
rect 23233 35332 23237 35388
rect 23173 35328 23237 35332
rect 23253 35388 23317 35392
rect 23253 35332 23257 35388
rect 23257 35332 23313 35388
rect 23313 35332 23317 35388
rect 23253 35328 23317 35332
rect 23333 35388 23397 35392
rect 23333 35332 23337 35388
rect 23337 35332 23393 35388
rect 23393 35332 23397 35388
rect 23333 35328 23397 35332
rect 6487 34844 6551 34848
rect 6487 34788 6491 34844
rect 6491 34788 6547 34844
rect 6547 34788 6551 34844
rect 6487 34784 6551 34788
rect 6567 34844 6631 34848
rect 6567 34788 6571 34844
rect 6571 34788 6627 34844
rect 6627 34788 6631 34844
rect 6567 34784 6631 34788
rect 6647 34844 6711 34848
rect 6647 34788 6651 34844
rect 6651 34788 6707 34844
rect 6707 34788 6711 34844
rect 6647 34784 6711 34788
rect 6727 34844 6791 34848
rect 6727 34788 6731 34844
rect 6731 34788 6787 34844
rect 6787 34788 6791 34844
rect 6727 34784 6791 34788
rect 17558 34844 17622 34848
rect 17558 34788 17562 34844
rect 17562 34788 17618 34844
rect 17618 34788 17622 34844
rect 17558 34784 17622 34788
rect 17638 34844 17702 34848
rect 17638 34788 17642 34844
rect 17642 34788 17698 34844
rect 17698 34788 17702 34844
rect 17638 34784 17702 34788
rect 17718 34844 17782 34848
rect 17718 34788 17722 34844
rect 17722 34788 17778 34844
rect 17778 34788 17782 34844
rect 17718 34784 17782 34788
rect 17798 34844 17862 34848
rect 17798 34788 17802 34844
rect 17802 34788 17858 34844
rect 17858 34788 17862 34844
rect 17798 34784 17862 34788
rect 28628 34844 28692 34848
rect 28628 34788 28632 34844
rect 28632 34788 28688 34844
rect 28688 34788 28692 34844
rect 28628 34784 28692 34788
rect 28708 34844 28772 34848
rect 28708 34788 28712 34844
rect 28712 34788 28768 34844
rect 28768 34788 28772 34844
rect 28708 34784 28772 34788
rect 28788 34844 28852 34848
rect 28788 34788 28792 34844
rect 28792 34788 28848 34844
rect 28848 34788 28852 34844
rect 28788 34784 28852 34788
rect 28868 34844 28932 34848
rect 28868 34788 28872 34844
rect 28872 34788 28928 34844
rect 28928 34788 28932 34844
rect 28868 34784 28932 34788
rect 12022 34300 12086 34304
rect 12022 34244 12026 34300
rect 12026 34244 12082 34300
rect 12082 34244 12086 34300
rect 12022 34240 12086 34244
rect 12102 34300 12166 34304
rect 12102 34244 12106 34300
rect 12106 34244 12162 34300
rect 12162 34244 12166 34300
rect 12102 34240 12166 34244
rect 12182 34300 12246 34304
rect 12182 34244 12186 34300
rect 12186 34244 12242 34300
rect 12242 34244 12246 34300
rect 12182 34240 12246 34244
rect 12262 34300 12326 34304
rect 12262 34244 12266 34300
rect 12266 34244 12322 34300
rect 12322 34244 12326 34300
rect 12262 34240 12326 34244
rect 23093 34300 23157 34304
rect 23093 34244 23097 34300
rect 23097 34244 23153 34300
rect 23153 34244 23157 34300
rect 23093 34240 23157 34244
rect 23173 34300 23237 34304
rect 23173 34244 23177 34300
rect 23177 34244 23233 34300
rect 23233 34244 23237 34300
rect 23173 34240 23237 34244
rect 23253 34300 23317 34304
rect 23253 34244 23257 34300
rect 23257 34244 23313 34300
rect 23313 34244 23317 34300
rect 23253 34240 23317 34244
rect 23333 34300 23397 34304
rect 23333 34244 23337 34300
rect 23337 34244 23393 34300
rect 23393 34244 23397 34300
rect 23333 34240 23397 34244
rect 6487 33756 6551 33760
rect 6487 33700 6491 33756
rect 6491 33700 6547 33756
rect 6547 33700 6551 33756
rect 6487 33696 6551 33700
rect 6567 33756 6631 33760
rect 6567 33700 6571 33756
rect 6571 33700 6627 33756
rect 6627 33700 6631 33756
rect 6567 33696 6631 33700
rect 6647 33756 6711 33760
rect 6647 33700 6651 33756
rect 6651 33700 6707 33756
rect 6707 33700 6711 33756
rect 6647 33696 6711 33700
rect 6727 33756 6791 33760
rect 6727 33700 6731 33756
rect 6731 33700 6787 33756
rect 6787 33700 6791 33756
rect 6727 33696 6791 33700
rect 17558 33756 17622 33760
rect 17558 33700 17562 33756
rect 17562 33700 17618 33756
rect 17618 33700 17622 33756
rect 17558 33696 17622 33700
rect 17638 33756 17702 33760
rect 17638 33700 17642 33756
rect 17642 33700 17698 33756
rect 17698 33700 17702 33756
rect 17638 33696 17702 33700
rect 17718 33756 17782 33760
rect 17718 33700 17722 33756
rect 17722 33700 17778 33756
rect 17778 33700 17782 33756
rect 17718 33696 17782 33700
rect 17798 33756 17862 33760
rect 17798 33700 17802 33756
rect 17802 33700 17858 33756
rect 17858 33700 17862 33756
rect 17798 33696 17862 33700
rect 28628 33756 28692 33760
rect 28628 33700 28632 33756
rect 28632 33700 28688 33756
rect 28688 33700 28692 33756
rect 28628 33696 28692 33700
rect 28708 33756 28772 33760
rect 28708 33700 28712 33756
rect 28712 33700 28768 33756
rect 28768 33700 28772 33756
rect 28708 33696 28772 33700
rect 28788 33756 28852 33760
rect 28788 33700 28792 33756
rect 28792 33700 28848 33756
rect 28848 33700 28852 33756
rect 28788 33696 28852 33700
rect 28868 33756 28932 33760
rect 28868 33700 28872 33756
rect 28872 33700 28928 33756
rect 28928 33700 28932 33756
rect 28868 33696 28932 33700
rect 12022 33212 12086 33216
rect 12022 33156 12026 33212
rect 12026 33156 12082 33212
rect 12082 33156 12086 33212
rect 12022 33152 12086 33156
rect 12102 33212 12166 33216
rect 12102 33156 12106 33212
rect 12106 33156 12162 33212
rect 12162 33156 12166 33212
rect 12102 33152 12166 33156
rect 12182 33212 12246 33216
rect 12182 33156 12186 33212
rect 12186 33156 12242 33212
rect 12242 33156 12246 33212
rect 12182 33152 12246 33156
rect 12262 33212 12326 33216
rect 12262 33156 12266 33212
rect 12266 33156 12322 33212
rect 12322 33156 12326 33212
rect 12262 33152 12326 33156
rect 23093 33212 23157 33216
rect 23093 33156 23097 33212
rect 23097 33156 23153 33212
rect 23153 33156 23157 33212
rect 23093 33152 23157 33156
rect 23173 33212 23237 33216
rect 23173 33156 23177 33212
rect 23177 33156 23233 33212
rect 23233 33156 23237 33212
rect 23173 33152 23237 33156
rect 23253 33212 23317 33216
rect 23253 33156 23257 33212
rect 23257 33156 23313 33212
rect 23313 33156 23317 33212
rect 23253 33152 23317 33156
rect 23333 33212 23397 33216
rect 23333 33156 23337 33212
rect 23337 33156 23393 33212
rect 23393 33156 23397 33212
rect 23333 33152 23397 33156
rect 6487 32668 6551 32672
rect 6487 32612 6491 32668
rect 6491 32612 6547 32668
rect 6547 32612 6551 32668
rect 6487 32608 6551 32612
rect 6567 32668 6631 32672
rect 6567 32612 6571 32668
rect 6571 32612 6627 32668
rect 6627 32612 6631 32668
rect 6567 32608 6631 32612
rect 6647 32668 6711 32672
rect 6647 32612 6651 32668
rect 6651 32612 6707 32668
rect 6707 32612 6711 32668
rect 6647 32608 6711 32612
rect 6727 32668 6791 32672
rect 6727 32612 6731 32668
rect 6731 32612 6787 32668
rect 6787 32612 6791 32668
rect 6727 32608 6791 32612
rect 17558 32668 17622 32672
rect 17558 32612 17562 32668
rect 17562 32612 17618 32668
rect 17618 32612 17622 32668
rect 17558 32608 17622 32612
rect 17638 32668 17702 32672
rect 17638 32612 17642 32668
rect 17642 32612 17698 32668
rect 17698 32612 17702 32668
rect 17638 32608 17702 32612
rect 17718 32668 17782 32672
rect 17718 32612 17722 32668
rect 17722 32612 17778 32668
rect 17778 32612 17782 32668
rect 17718 32608 17782 32612
rect 17798 32668 17862 32672
rect 17798 32612 17802 32668
rect 17802 32612 17858 32668
rect 17858 32612 17862 32668
rect 17798 32608 17862 32612
rect 28628 32668 28692 32672
rect 28628 32612 28632 32668
rect 28632 32612 28688 32668
rect 28688 32612 28692 32668
rect 28628 32608 28692 32612
rect 28708 32668 28772 32672
rect 28708 32612 28712 32668
rect 28712 32612 28768 32668
rect 28768 32612 28772 32668
rect 28708 32608 28772 32612
rect 28788 32668 28852 32672
rect 28788 32612 28792 32668
rect 28792 32612 28848 32668
rect 28848 32612 28852 32668
rect 28788 32608 28852 32612
rect 28868 32668 28932 32672
rect 28868 32612 28872 32668
rect 28872 32612 28928 32668
rect 28928 32612 28932 32668
rect 28868 32608 28932 32612
rect 12022 32124 12086 32128
rect 12022 32068 12026 32124
rect 12026 32068 12082 32124
rect 12082 32068 12086 32124
rect 12022 32064 12086 32068
rect 12102 32124 12166 32128
rect 12102 32068 12106 32124
rect 12106 32068 12162 32124
rect 12162 32068 12166 32124
rect 12102 32064 12166 32068
rect 12182 32124 12246 32128
rect 12182 32068 12186 32124
rect 12186 32068 12242 32124
rect 12242 32068 12246 32124
rect 12182 32064 12246 32068
rect 12262 32124 12326 32128
rect 12262 32068 12266 32124
rect 12266 32068 12322 32124
rect 12322 32068 12326 32124
rect 12262 32064 12326 32068
rect 23093 32124 23157 32128
rect 23093 32068 23097 32124
rect 23097 32068 23153 32124
rect 23153 32068 23157 32124
rect 23093 32064 23157 32068
rect 23173 32124 23237 32128
rect 23173 32068 23177 32124
rect 23177 32068 23233 32124
rect 23233 32068 23237 32124
rect 23173 32064 23237 32068
rect 23253 32124 23317 32128
rect 23253 32068 23257 32124
rect 23257 32068 23313 32124
rect 23313 32068 23317 32124
rect 23253 32064 23317 32068
rect 23333 32124 23397 32128
rect 23333 32068 23337 32124
rect 23337 32068 23393 32124
rect 23393 32068 23397 32124
rect 23333 32064 23397 32068
rect 6487 31580 6551 31584
rect 6487 31524 6491 31580
rect 6491 31524 6547 31580
rect 6547 31524 6551 31580
rect 6487 31520 6551 31524
rect 6567 31580 6631 31584
rect 6567 31524 6571 31580
rect 6571 31524 6627 31580
rect 6627 31524 6631 31580
rect 6567 31520 6631 31524
rect 6647 31580 6711 31584
rect 6647 31524 6651 31580
rect 6651 31524 6707 31580
rect 6707 31524 6711 31580
rect 6647 31520 6711 31524
rect 6727 31580 6791 31584
rect 6727 31524 6731 31580
rect 6731 31524 6787 31580
rect 6787 31524 6791 31580
rect 6727 31520 6791 31524
rect 17558 31580 17622 31584
rect 17558 31524 17562 31580
rect 17562 31524 17618 31580
rect 17618 31524 17622 31580
rect 17558 31520 17622 31524
rect 17638 31580 17702 31584
rect 17638 31524 17642 31580
rect 17642 31524 17698 31580
rect 17698 31524 17702 31580
rect 17638 31520 17702 31524
rect 17718 31580 17782 31584
rect 17718 31524 17722 31580
rect 17722 31524 17778 31580
rect 17778 31524 17782 31580
rect 17718 31520 17782 31524
rect 17798 31580 17862 31584
rect 17798 31524 17802 31580
rect 17802 31524 17858 31580
rect 17858 31524 17862 31580
rect 17798 31520 17862 31524
rect 28628 31580 28692 31584
rect 28628 31524 28632 31580
rect 28632 31524 28688 31580
rect 28688 31524 28692 31580
rect 28628 31520 28692 31524
rect 28708 31580 28772 31584
rect 28708 31524 28712 31580
rect 28712 31524 28768 31580
rect 28768 31524 28772 31580
rect 28708 31520 28772 31524
rect 28788 31580 28852 31584
rect 28788 31524 28792 31580
rect 28792 31524 28848 31580
rect 28848 31524 28852 31580
rect 28788 31520 28852 31524
rect 28868 31580 28932 31584
rect 28868 31524 28872 31580
rect 28872 31524 28928 31580
rect 28928 31524 28932 31580
rect 28868 31520 28932 31524
rect 12022 31036 12086 31040
rect 12022 30980 12026 31036
rect 12026 30980 12082 31036
rect 12082 30980 12086 31036
rect 12022 30976 12086 30980
rect 12102 31036 12166 31040
rect 12102 30980 12106 31036
rect 12106 30980 12162 31036
rect 12162 30980 12166 31036
rect 12102 30976 12166 30980
rect 12182 31036 12246 31040
rect 12182 30980 12186 31036
rect 12186 30980 12242 31036
rect 12242 30980 12246 31036
rect 12182 30976 12246 30980
rect 12262 31036 12326 31040
rect 12262 30980 12266 31036
rect 12266 30980 12322 31036
rect 12322 30980 12326 31036
rect 12262 30976 12326 30980
rect 23093 31036 23157 31040
rect 23093 30980 23097 31036
rect 23097 30980 23153 31036
rect 23153 30980 23157 31036
rect 23093 30976 23157 30980
rect 23173 31036 23237 31040
rect 23173 30980 23177 31036
rect 23177 30980 23233 31036
rect 23233 30980 23237 31036
rect 23173 30976 23237 30980
rect 23253 31036 23317 31040
rect 23253 30980 23257 31036
rect 23257 30980 23313 31036
rect 23313 30980 23317 31036
rect 23253 30976 23317 30980
rect 23333 31036 23397 31040
rect 23333 30980 23337 31036
rect 23337 30980 23393 31036
rect 23393 30980 23397 31036
rect 23333 30976 23397 30980
rect 6487 30492 6551 30496
rect 6487 30436 6491 30492
rect 6491 30436 6547 30492
rect 6547 30436 6551 30492
rect 6487 30432 6551 30436
rect 6567 30492 6631 30496
rect 6567 30436 6571 30492
rect 6571 30436 6627 30492
rect 6627 30436 6631 30492
rect 6567 30432 6631 30436
rect 6647 30492 6711 30496
rect 6647 30436 6651 30492
rect 6651 30436 6707 30492
rect 6707 30436 6711 30492
rect 6647 30432 6711 30436
rect 6727 30492 6791 30496
rect 6727 30436 6731 30492
rect 6731 30436 6787 30492
rect 6787 30436 6791 30492
rect 6727 30432 6791 30436
rect 17558 30492 17622 30496
rect 17558 30436 17562 30492
rect 17562 30436 17618 30492
rect 17618 30436 17622 30492
rect 17558 30432 17622 30436
rect 17638 30492 17702 30496
rect 17638 30436 17642 30492
rect 17642 30436 17698 30492
rect 17698 30436 17702 30492
rect 17638 30432 17702 30436
rect 17718 30492 17782 30496
rect 17718 30436 17722 30492
rect 17722 30436 17778 30492
rect 17778 30436 17782 30492
rect 17718 30432 17782 30436
rect 17798 30492 17862 30496
rect 17798 30436 17802 30492
rect 17802 30436 17858 30492
rect 17858 30436 17862 30492
rect 17798 30432 17862 30436
rect 28628 30492 28692 30496
rect 28628 30436 28632 30492
rect 28632 30436 28688 30492
rect 28688 30436 28692 30492
rect 28628 30432 28692 30436
rect 28708 30492 28772 30496
rect 28708 30436 28712 30492
rect 28712 30436 28768 30492
rect 28768 30436 28772 30492
rect 28708 30432 28772 30436
rect 28788 30492 28852 30496
rect 28788 30436 28792 30492
rect 28792 30436 28848 30492
rect 28848 30436 28852 30492
rect 28788 30432 28852 30436
rect 28868 30492 28932 30496
rect 28868 30436 28872 30492
rect 28872 30436 28928 30492
rect 28928 30436 28932 30492
rect 28868 30432 28932 30436
rect 12022 29948 12086 29952
rect 12022 29892 12026 29948
rect 12026 29892 12082 29948
rect 12082 29892 12086 29948
rect 12022 29888 12086 29892
rect 12102 29948 12166 29952
rect 12102 29892 12106 29948
rect 12106 29892 12162 29948
rect 12162 29892 12166 29948
rect 12102 29888 12166 29892
rect 12182 29948 12246 29952
rect 12182 29892 12186 29948
rect 12186 29892 12242 29948
rect 12242 29892 12246 29948
rect 12182 29888 12246 29892
rect 12262 29948 12326 29952
rect 12262 29892 12266 29948
rect 12266 29892 12322 29948
rect 12322 29892 12326 29948
rect 12262 29888 12326 29892
rect 23093 29948 23157 29952
rect 23093 29892 23097 29948
rect 23097 29892 23153 29948
rect 23153 29892 23157 29948
rect 23093 29888 23157 29892
rect 23173 29948 23237 29952
rect 23173 29892 23177 29948
rect 23177 29892 23233 29948
rect 23233 29892 23237 29948
rect 23173 29888 23237 29892
rect 23253 29948 23317 29952
rect 23253 29892 23257 29948
rect 23257 29892 23313 29948
rect 23313 29892 23317 29948
rect 23253 29888 23317 29892
rect 23333 29948 23397 29952
rect 23333 29892 23337 29948
rect 23337 29892 23393 29948
rect 23393 29892 23397 29948
rect 23333 29888 23397 29892
rect 6487 29404 6551 29408
rect 6487 29348 6491 29404
rect 6491 29348 6547 29404
rect 6547 29348 6551 29404
rect 6487 29344 6551 29348
rect 6567 29404 6631 29408
rect 6567 29348 6571 29404
rect 6571 29348 6627 29404
rect 6627 29348 6631 29404
rect 6567 29344 6631 29348
rect 6647 29404 6711 29408
rect 6647 29348 6651 29404
rect 6651 29348 6707 29404
rect 6707 29348 6711 29404
rect 6647 29344 6711 29348
rect 6727 29404 6791 29408
rect 6727 29348 6731 29404
rect 6731 29348 6787 29404
rect 6787 29348 6791 29404
rect 6727 29344 6791 29348
rect 17558 29404 17622 29408
rect 17558 29348 17562 29404
rect 17562 29348 17618 29404
rect 17618 29348 17622 29404
rect 17558 29344 17622 29348
rect 17638 29404 17702 29408
rect 17638 29348 17642 29404
rect 17642 29348 17698 29404
rect 17698 29348 17702 29404
rect 17638 29344 17702 29348
rect 17718 29404 17782 29408
rect 17718 29348 17722 29404
rect 17722 29348 17778 29404
rect 17778 29348 17782 29404
rect 17718 29344 17782 29348
rect 17798 29404 17862 29408
rect 17798 29348 17802 29404
rect 17802 29348 17858 29404
rect 17858 29348 17862 29404
rect 17798 29344 17862 29348
rect 28628 29404 28692 29408
rect 28628 29348 28632 29404
rect 28632 29348 28688 29404
rect 28688 29348 28692 29404
rect 28628 29344 28692 29348
rect 28708 29404 28772 29408
rect 28708 29348 28712 29404
rect 28712 29348 28768 29404
rect 28768 29348 28772 29404
rect 28708 29344 28772 29348
rect 28788 29404 28852 29408
rect 28788 29348 28792 29404
rect 28792 29348 28848 29404
rect 28848 29348 28852 29404
rect 28788 29344 28852 29348
rect 28868 29404 28932 29408
rect 28868 29348 28872 29404
rect 28872 29348 28928 29404
rect 28928 29348 28932 29404
rect 28868 29344 28932 29348
rect 12022 28860 12086 28864
rect 12022 28804 12026 28860
rect 12026 28804 12082 28860
rect 12082 28804 12086 28860
rect 12022 28800 12086 28804
rect 12102 28860 12166 28864
rect 12102 28804 12106 28860
rect 12106 28804 12162 28860
rect 12162 28804 12166 28860
rect 12102 28800 12166 28804
rect 12182 28860 12246 28864
rect 12182 28804 12186 28860
rect 12186 28804 12242 28860
rect 12242 28804 12246 28860
rect 12182 28800 12246 28804
rect 12262 28860 12326 28864
rect 12262 28804 12266 28860
rect 12266 28804 12322 28860
rect 12322 28804 12326 28860
rect 12262 28800 12326 28804
rect 23093 28860 23157 28864
rect 23093 28804 23097 28860
rect 23097 28804 23153 28860
rect 23153 28804 23157 28860
rect 23093 28800 23157 28804
rect 23173 28860 23237 28864
rect 23173 28804 23177 28860
rect 23177 28804 23233 28860
rect 23233 28804 23237 28860
rect 23173 28800 23237 28804
rect 23253 28860 23317 28864
rect 23253 28804 23257 28860
rect 23257 28804 23313 28860
rect 23313 28804 23317 28860
rect 23253 28800 23317 28804
rect 23333 28860 23397 28864
rect 23333 28804 23337 28860
rect 23337 28804 23393 28860
rect 23393 28804 23397 28860
rect 23333 28800 23397 28804
rect 6487 28316 6551 28320
rect 6487 28260 6491 28316
rect 6491 28260 6547 28316
rect 6547 28260 6551 28316
rect 6487 28256 6551 28260
rect 6567 28316 6631 28320
rect 6567 28260 6571 28316
rect 6571 28260 6627 28316
rect 6627 28260 6631 28316
rect 6567 28256 6631 28260
rect 6647 28316 6711 28320
rect 6647 28260 6651 28316
rect 6651 28260 6707 28316
rect 6707 28260 6711 28316
rect 6647 28256 6711 28260
rect 6727 28316 6791 28320
rect 6727 28260 6731 28316
rect 6731 28260 6787 28316
rect 6787 28260 6791 28316
rect 6727 28256 6791 28260
rect 17558 28316 17622 28320
rect 17558 28260 17562 28316
rect 17562 28260 17618 28316
rect 17618 28260 17622 28316
rect 17558 28256 17622 28260
rect 17638 28316 17702 28320
rect 17638 28260 17642 28316
rect 17642 28260 17698 28316
rect 17698 28260 17702 28316
rect 17638 28256 17702 28260
rect 17718 28316 17782 28320
rect 17718 28260 17722 28316
rect 17722 28260 17778 28316
rect 17778 28260 17782 28316
rect 17718 28256 17782 28260
rect 17798 28316 17862 28320
rect 17798 28260 17802 28316
rect 17802 28260 17858 28316
rect 17858 28260 17862 28316
rect 17798 28256 17862 28260
rect 28628 28316 28692 28320
rect 28628 28260 28632 28316
rect 28632 28260 28688 28316
rect 28688 28260 28692 28316
rect 28628 28256 28692 28260
rect 28708 28316 28772 28320
rect 28708 28260 28712 28316
rect 28712 28260 28768 28316
rect 28768 28260 28772 28316
rect 28708 28256 28772 28260
rect 28788 28316 28852 28320
rect 28788 28260 28792 28316
rect 28792 28260 28848 28316
rect 28848 28260 28852 28316
rect 28788 28256 28852 28260
rect 28868 28316 28932 28320
rect 28868 28260 28872 28316
rect 28872 28260 28928 28316
rect 28928 28260 28932 28316
rect 28868 28256 28932 28260
rect 12022 27772 12086 27776
rect 12022 27716 12026 27772
rect 12026 27716 12082 27772
rect 12082 27716 12086 27772
rect 12022 27712 12086 27716
rect 12102 27772 12166 27776
rect 12102 27716 12106 27772
rect 12106 27716 12162 27772
rect 12162 27716 12166 27772
rect 12102 27712 12166 27716
rect 12182 27772 12246 27776
rect 12182 27716 12186 27772
rect 12186 27716 12242 27772
rect 12242 27716 12246 27772
rect 12182 27712 12246 27716
rect 12262 27772 12326 27776
rect 12262 27716 12266 27772
rect 12266 27716 12322 27772
rect 12322 27716 12326 27772
rect 12262 27712 12326 27716
rect 23093 27772 23157 27776
rect 23093 27716 23097 27772
rect 23097 27716 23153 27772
rect 23153 27716 23157 27772
rect 23093 27712 23157 27716
rect 23173 27772 23237 27776
rect 23173 27716 23177 27772
rect 23177 27716 23233 27772
rect 23233 27716 23237 27772
rect 23173 27712 23237 27716
rect 23253 27772 23317 27776
rect 23253 27716 23257 27772
rect 23257 27716 23313 27772
rect 23313 27716 23317 27772
rect 23253 27712 23317 27716
rect 23333 27772 23397 27776
rect 23333 27716 23337 27772
rect 23337 27716 23393 27772
rect 23393 27716 23397 27772
rect 23333 27712 23397 27716
rect 6487 27228 6551 27232
rect 6487 27172 6491 27228
rect 6491 27172 6547 27228
rect 6547 27172 6551 27228
rect 6487 27168 6551 27172
rect 6567 27228 6631 27232
rect 6567 27172 6571 27228
rect 6571 27172 6627 27228
rect 6627 27172 6631 27228
rect 6567 27168 6631 27172
rect 6647 27228 6711 27232
rect 6647 27172 6651 27228
rect 6651 27172 6707 27228
rect 6707 27172 6711 27228
rect 6647 27168 6711 27172
rect 6727 27228 6791 27232
rect 6727 27172 6731 27228
rect 6731 27172 6787 27228
rect 6787 27172 6791 27228
rect 6727 27168 6791 27172
rect 17558 27228 17622 27232
rect 17558 27172 17562 27228
rect 17562 27172 17618 27228
rect 17618 27172 17622 27228
rect 17558 27168 17622 27172
rect 17638 27228 17702 27232
rect 17638 27172 17642 27228
rect 17642 27172 17698 27228
rect 17698 27172 17702 27228
rect 17638 27168 17702 27172
rect 17718 27228 17782 27232
rect 17718 27172 17722 27228
rect 17722 27172 17778 27228
rect 17778 27172 17782 27228
rect 17718 27168 17782 27172
rect 17798 27228 17862 27232
rect 17798 27172 17802 27228
rect 17802 27172 17858 27228
rect 17858 27172 17862 27228
rect 17798 27168 17862 27172
rect 28628 27228 28692 27232
rect 28628 27172 28632 27228
rect 28632 27172 28688 27228
rect 28688 27172 28692 27228
rect 28628 27168 28692 27172
rect 28708 27228 28772 27232
rect 28708 27172 28712 27228
rect 28712 27172 28768 27228
rect 28768 27172 28772 27228
rect 28708 27168 28772 27172
rect 28788 27228 28852 27232
rect 28788 27172 28792 27228
rect 28792 27172 28848 27228
rect 28848 27172 28852 27228
rect 28788 27168 28852 27172
rect 28868 27228 28932 27232
rect 28868 27172 28872 27228
rect 28872 27172 28928 27228
rect 28928 27172 28932 27228
rect 28868 27168 28932 27172
rect 12022 26684 12086 26688
rect 12022 26628 12026 26684
rect 12026 26628 12082 26684
rect 12082 26628 12086 26684
rect 12022 26624 12086 26628
rect 12102 26684 12166 26688
rect 12102 26628 12106 26684
rect 12106 26628 12162 26684
rect 12162 26628 12166 26684
rect 12102 26624 12166 26628
rect 12182 26684 12246 26688
rect 12182 26628 12186 26684
rect 12186 26628 12242 26684
rect 12242 26628 12246 26684
rect 12182 26624 12246 26628
rect 12262 26684 12326 26688
rect 12262 26628 12266 26684
rect 12266 26628 12322 26684
rect 12322 26628 12326 26684
rect 12262 26624 12326 26628
rect 23093 26684 23157 26688
rect 23093 26628 23097 26684
rect 23097 26628 23153 26684
rect 23153 26628 23157 26684
rect 23093 26624 23157 26628
rect 23173 26684 23237 26688
rect 23173 26628 23177 26684
rect 23177 26628 23233 26684
rect 23233 26628 23237 26684
rect 23173 26624 23237 26628
rect 23253 26684 23317 26688
rect 23253 26628 23257 26684
rect 23257 26628 23313 26684
rect 23313 26628 23317 26684
rect 23253 26624 23317 26628
rect 23333 26684 23397 26688
rect 23333 26628 23337 26684
rect 23337 26628 23393 26684
rect 23393 26628 23397 26684
rect 23333 26624 23397 26628
rect 6487 26140 6551 26144
rect 6487 26084 6491 26140
rect 6491 26084 6547 26140
rect 6547 26084 6551 26140
rect 6487 26080 6551 26084
rect 6567 26140 6631 26144
rect 6567 26084 6571 26140
rect 6571 26084 6627 26140
rect 6627 26084 6631 26140
rect 6567 26080 6631 26084
rect 6647 26140 6711 26144
rect 6647 26084 6651 26140
rect 6651 26084 6707 26140
rect 6707 26084 6711 26140
rect 6647 26080 6711 26084
rect 6727 26140 6791 26144
rect 6727 26084 6731 26140
rect 6731 26084 6787 26140
rect 6787 26084 6791 26140
rect 6727 26080 6791 26084
rect 17558 26140 17622 26144
rect 17558 26084 17562 26140
rect 17562 26084 17618 26140
rect 17618 26084 17622 26140
rect 17558 26080 17622 26084
rect 17638 26140 17702 26144
rect 17638 26084 17642 26140
rect 17642 26084 17698 26140
rect 17698 26084 17702 26140
rect 17638 26080 17702 26084
rect 17718 26140 17782 26144
rect 17718 26084 17722 26140
rect 17722 26084 17778 26140
rect 17778 26084 17782 26140
rect 17718 26080 17782 26084
rect 17798 26140 17862 26144
rect 17798 26084 17802 26140
rect 17802 26084 17858 26140
rect 17858 26084 17862 26140
rect 17798 26080 17862 26084
rect 28628 26140 28692 26144
rect 28628 26084 28632 26140
rect 28632 26084 28688 26140
rect 28688 26084 28692 26140
rect 28628 26080 28692 26084
rect 28708 26140 28772 26144
rect 28708 26084 28712 26140
rect 28712 26084 28768 26140
rect 28768 26084 28772 26140
rect 28708 26080 28772 26084
rect 28788 26140 28852 26144
rect 28788 26084 28792 26140
rect 28792 26084 28848 26140
rect 28848 26084 28852 26140
rect 28788 26080 28852 26084
rect 28868 26140 28932 26144
rect 28868 26084 28872 26140
rect 28872 26084 28928 26140
rect 28928 26084 28932 26140
rect 28868 26080 28932 26084
rect 12022 25596 12086 25600
rect 12022 25540 12026 25596
rect 12026 25540 12082 25596
rect 12082 25540 12086 25596
rect 12022 25536 12086 25540
rect 12102 25596 12166 25600
rect 12102 25540 12106 25596
rect 12106 25540 12162 25596
rect 12162 25540 12166 25596
rect 12102 25536 12166 25540
rect 12182 25596 12246 25600
rect 12182 25540 12186 25596
rect 12186 25540 12242 25596
rect 12242 25540 12246 25596
rect 12182 25536 12246 25540
rect 12262 25596 12326 25600
rect 12262 25540 12266 25596
rect 12266 25540 12322 25596
rect 12322 25540 12326 25596
rect 12262 25536 12326 25540
rect 23093 25596 23157 25600
rect 23093 25540 23097 25596
rect 23097 25540 23153 25596
rect 23153 25540 23157 25596
rect 23093 25536 23157 25540
rect 23173 25596 23237 25600
rect 23173 25540 23177 25596
rect 23177 25540 23233 25596
rect 23233 25540 23237 25596
rect 23173 25536 23237 25540
rect 23253 25596 23317 25600
rect 23253 25540 23257 25596
rect 23257 25540 23313 25596
rect 23313 25540 23317 25596
rect 23253 25536 23317 25540
rect 23333 25596 23397 25600
rect 23333 25540 23337 25596
rect 23337 25540 23393 25596
rect 23393 25540 23397 25596
rect 23333 25536 23397 25540
rect 6487 25052 6551 25056
rect 6487 24996 6491 25052
rect 6491 24996 6547 25052
rect 6547 24996 6551 25052
rect 6487 24992 6551 24996
rect 6567 25052 6631 25056
rect 6567 24996 6571 25052
rect 6571 24996 6627 25052
rect 6627 24996 6631 25052
rect 6567 24992 6631 24996
rect 6647 25052 6711 25056
rect 6647 24996 6651 25052
rect 6651 24996 6707 25052
rect 6707 24996 6711 25052
rect 6647 24992 6711 24996
rect 6727 25052 6791 25056
rect 6727 24996 6731 25052
rect 6731 24996 6787 25052
rect 6787 24996 6791 25052
rect 6727 24992 6791 24996
rect 17558 25052 17622 25056
rect 17558 24996 17562 25052
rect 17562 24996 17618 25052
rect 17618 24996 17622 25052
rect 17558 24992 17622 24996
rect 17638 25052 17702 25056
rect 17638 24996 17642 25052
rect 17642 24996 17698 25052
rect 17698 24996 17702 25052
rect 17638 24992 17702 24996
rect 17718 25052 17782 25056
rect 17718 24996 17722 25052
rect 17722 24996 17778 25052
rect 17778 24996 17782 25052
rect 17718 24992 17782 24996
rect 17798 25052 17862 25056
rect 17798 24996 17802 25052
rect 17802 24996 17858 25052
rect 17858 24996 17862 25052
rect 17798 24992 17862 24996
rect 28628 25052 28692 25056
rect 28628 24996 28632 25052
rect 28632 24996 28688 25052
rect 28688 24996 28692 25052
rect 28628 24992 28692 24996
rect 28708 25052 28772 25056
rect 28708 24996 28712 25052
rect 28712 24996 28768 25052
rect 28768 24996 28772 25052
rect 28708 24992 28772 24996
rect 28788 25052 28852 25056
rect 28788 24996 28792 25052
rect 28792 24996 28848 25052
rect 28848 24996 28852 25052
rect 28788 24992 28852 24996
rect 28868 25052 28932 25056
rect 28868 24996 28872 25052
rect 28872 24996 28928 25052
rect 28928 24996 28932 25052
rect 28868 24992 28932 24996
rect 12022 24508 12086 24512
rect 12022 24452 12026 24508
rect 12026 24452 12082 24508
rect 12082 24452 12086 24508
rect 12022 24448 12086 24452
rect 12102 24508 12166 24512
rect 12102 24452 12106 24508
rect 12106 24452 12162 24508
rect 12162 24452 12166 24508
rect 12102 24448 12166 24452
rect 12182 24508 12246 24512
rect 12182 24452 12186 24508
rect 12186 24452 12242 24508
rect 12242 24452 12246 24508
rect 12182 24448 12246 24452
rect 12262 24508 12326 24512
rect 12262 24452 12266 24508
rect 12266 24452 12322 24508
rect 12322 24452 12326 24508
rect 12262 24448 12326 24452
rect 23093 24508 23157 24512
rect 23093 24452 23097 24508
rect 23097 24452 23153 24508
rect 23153 24452 23157 24508
rect 23093 24448 23157 24452
rect 23173 24508 23237 24512
rect 23173 24452 23177 24508
rect 23177 24452 23233 24508
rect 23233 24452 23237 24508
rect 23173 24448 23237 24452
rect 23253 24508 23317 24512
rect 23253 24452 23257 24508
rect 23257 24452 23313 24508
rect 23313 24452 23317 24508
rect 23253 24448 23317 24452
rect 23333 24508 23397 24512
rect 23333 24452 23337 24508
rect 23337 24452 23393 24508
rect 23393 24452 23397 24508
rect 23333 24448 23397 24452
rect 6487 23964 6551 23968
rect 6487 23908 6491 23964
rect 6491 23908 6547 23964
rect 6547 23908 6551 23964
rect 6487 23904 6551 23908
rect 6567 23964 6631 23968
rect 6567 23908 6571 23964
rect 6571 23908 6627 23964
rect 6627 23908 6631 23964
rect 6567 23904 6631 23908
rect 6647 23964 6711 23968
rect 6647 23908 6651 23964
rect 6651 23908 6707 23964
rect 6707 23908 6711 23964
rect 6647 23904 6711 23908
rect 6727 23964 6791 23968
rect 6727 23908 6731 23964
rect 6731 23908 6787 23964
rect 6787 23908 6791 23964
rect 6727 23904 6791 23908
rect 17558 23964 17622 23968
rect 17558 23908 17562 23964
rect 17562 23908 17618 23964
rect 17618 23908 17622 23964
rect 17558 23904 17622 23908
rect 17638 23964 17702 23968
rect 17638 23908 17642 23964
rect 17642 23908 17698 23964
rect 17698 23908 17702 23964
rect 17638 23904 17702 23908
rect 17718 23964 17782 23968
rect 17718 23908 17722 23964
rect 17722 23908 17778 23964
rect 17778 23908 17782 23964
rect 17718 23904 17782 23908
rect 17798 23964 17862 23968
rect 17798 23908 17802 23964
rect 17802 23908 17858 23964
rect 17858 23908 17862 23964
rect 17798 23904 17862 23908
rect 28628 23964 28692 23968
rect 28628 23908 28632 23964
rect 28632 23908 28688 23964
rect 28688 23908 28692 23964
rect 28628 23904 28692 23908
rect 28708 23964 28772 23968
rect 28708 23908 28712 23964
rect 28712 23908 28768 23964
rect 28768 23908 28772 23964
rect 28708 23904 28772 23908
rect 28788 23964 28852 23968
rect 28788 23908 28792 23964
rect 28792 23908 28848 23964
rect 28848 23908 28852 23964
rect 28788 23904 28852 23908
rect 28868 23964 28932 23968
rect 28868 23908 28872 23964
rect 28872 23908 28928 23964
rect 28928 23908 28932 23964
rect 28868 23904 28932 23908
rect 12022 23420 12086 23424
rect 12022 23364 12026 23420
rect 12026 23364 12082 23420
rect 12082 23364 12086 23420
rect 12022 23360 12086 23364
rect 12102 23420 12166 23424
rect 12102 23364 12106 23420
rect 12106 23364 12162 23420
rect 12162 23364 12166 23420
rect 12102 23360 12166 23364
rect 12182 23420 12246 23424
rect 12182 23364 12186 23420
rect 12186 23364 12242 23420
rect 12242 23364 12246 23420
rect 12182 23360 12246 23364
rect 12262 23420 12326 23424
rect 12262 23364 12266 23420
rect 12266 23364 12322 23420
rect 12322 23364 12326 23420
rect 12262 23360 12326 23364
rect 23093 23420 23157 23424
rect 23093 23364 23097 23420
rect 23097 23364 23153 23420
rect 23153 23364 23157 23420
rect 23093 23360 23157 23364
rect 23173 23420 23237 23424
rect 23173 23364 23177 23420
rect 23177 23364 23233 23420
rect 23233 23364 23237 23420
rect 23173 23360 23237 23364
rect 23253 23420 23317 23424
rect 23253 23364 23257 23420
rect 23257 23364 23313 23420
rect 23313 23364 23317 23420
rect 23253 23360 23317 23364
rect 23333 23420 23397 23424
rect 23333 23364 23337 23420
rect 23337 23364 23393 23420
rect 23393 23364 23397 23420
rect 23333 23360 23397 23364
rect 6487 22876 6551 22880
rect 6487 22820 6491 22876
rect 6491 22820 6547 22876
rect 6547 22820 6551 22876
rect 6487 22816 6551 22820
rect 6567 22876 6631 22880
rect 6567 22820 6571 22876
rect 6571 22820 6627 22876
rect 6627 22820 6631 22876
rect 6567 22816 6631 22820
rect 6647 22876 6711 22880
rect 6647 22820 6651 22876
rect 6651 22820 6707 22876
rect 6707 22820 6711 22876
rect 6647 22816 6711 22820
rect 6727 22876 6791 22880
rect 6727 22820 6731 22876
rect 6731 22820 6787 22876
rect 6787 22820 6791 22876
rect 6727 22816 6791 22820
rect 17558 22876 17622 22880
rect 17558 22820 17562 22876
rect 17562 22820 17618 22876
rect 17618 22820 17622 22876
rect 17558 22816 17622 22820
rect 17638 22876 17702 22880
rect 17638 22820 17642 22876
rect 17642 22820 17698 22876
rect 17698 22820 17702 22876
rect 17638 22816 17702 22820
rect 17718 22876 17782 22880
rect 17718 22820 17722 22876
rect 17722 22820 17778 22876
rect 17778 22820 17782 22876
rect 17718 22816 17782 22820
rect 17798 22876 17862 22880
rect 17798 22820 17802 22876
rect 17802 22820 17858 22876
rect 17858 22820 17862 22876
rect 17798 22816 17862 22820
rect 28628 22876 28692 22880
rect 28628 22820 28632 22876
rect 28632 22820 28688 22876
rect 28688 22820 28692 22876
rect 28628 22816 28692 22820
rect 28708 22876 28772 22880
rect 28708 22820 28712 22876
rect 28712 22820 28768 22876
rect 28768 22820 28772 22876
rect 28708 22816 28772 22820
rect 28788 22876 28852 22880
rect 28788 22820 28792 22876
rect 28792 22820 28848 22876
rect 28848 22820 28852 22876
rect 28788 22816 28852 22820
rect 28868 22876 28932 22880
rect 28868 22820 28872 22876
rect 28872 22820 28928 22876
rect 28928 22820 28932 22876
rect 28868 22816 28932 22820
rect 12022 22332 12086 22336
rect 12022 22276 12026 22332
rect 12026 22276 12082 22332
rect 12082 22276 12086 22332
rect 12022 22272 12086 22276
rect 12102 22332 12166 22336
rect 12102 22276 12106 22332
rect 12106 22276 12162 22332
rect 12162 22276 12166 22332
rect 12102 22272 12166 22276
rect 12182 22332 12246 22336
rect 12182 22276 12186 22332
rect 12186 22276 12242 22332
rect 12242 22276 12246 22332
rect 12182 22272 12246 22276
rect 12262 22332 12326 22336
rect 12262 22276 12266 22332
rect 12266 22276 12322 22332
rect 12322 22276 12326 22332
rect 12262 22272 12326 22276
rect 23093 22332 23157 22336
rect 23093 22276 23097 22332
rect 23097 22276 23153 22332
rect 23153 22276 23157 22332
rect 23093 22272 23157 22276
rect 23173 22332 23237 22336
rect 23173 22276 23177 22332
rect 23177 22276 23233 22332
rect 23233 22276 23237 22332
rect 23173 22272 23237 22276
rect 23253 22332 23317 22336
rect 23253 22276 23257 22332
rect 23257 22276 23313 22332
rect 23313 22276 23317 22332
rect 23253 22272 23317 22276
rect 23333 22332 23397 22336
rect 23333 22276 23337 22332
rect 23337 22276 23393 22332
rect 23393 22276 23397 22332
rect 23333 22272 23397 22276
rect 6487 21788 6551 21792
rect 6487 21732 6491 21788
rect 6491 21732 6547 21788
rect 6547 21732 6551 21788
rect 6487 21728 6551 21732
rect 6567 21788 6631 21792
rect 6567 21732 6571 21788
rect 6571 21732 6627 21788
rect 6627 21732 6631 21788
rect 6567 21728 6631 21732
rect 6647 21788 6711 21792
rect 6647 21732 6651 21788
rect 6651 21732 6707 21788
rect 6707 21732 6711 21788
rect 6647 21728 6711 21732
rect 6727 21788 6791 21792
rect 6727 21732 6731 21788
rect 6731 21732 6787 21788
rect 6787 21732 6791 21788
rect 6727 21728 6791 21732
rect 17558 21788 17622 21792
rect 17558 21732 17562 21788
rect 17562 21732 17618 21788
rect 17618 21732 17622 21788
rect 17558 21728 17622 21732
rect 17638 21788 17702 21792
rect 17638 21732 17642 21788
rect 17642 21732 17698 21788
rect 17698 21732 17702 21788
rect 17638 21728 17702 21732
rect 17718 21788 17782 21792
rect 17718 21732 17722 21788
rect 17722 21732 17778 21788
rect 17778 21732 17782 21788
rect 17718 21728 17782 21732
rect 17798 21788 17862 21792
rect 17798 21732 17802 21788
rect 17802 21732 17858 21788
rect 17858 21732 17862 21788
rect 17798 21728 17862 21732
rect 28628 21788 28692 21792
rect 28628 21732 28632 21788
rect 28632 21732 28688 21788
rect 28688 21732 28692 21788
rect 28628 21728 28692 21732
rect 28708 21788 28772 21792
rect 28708 21732 28712 21788
rect 28712 21732 28768 21788
rect 28768 21732 28772 21788
rect 28708 21728 28772 21732
rect 28788 21788 28852 21792
rect 28788 21732 28792 21788
rect 28792 21732 28848 21788
rect 28848 21732 28852 21788
rect 28788 21728 28852 21732
rect 28868 21788 28932 21792
rect 28868 21732 28872 21788
rect 28872 21732 28928 21788
rect 28928 21732 28932 21788
rect 28868 21728 28932 21732
rect 12022 21244 12086 21248
rect 12022 21188 12026 21244
rect 12026 21188 12082 21244
rect 12082 21188 12086 21244
rect 12022 21184 12086 21188
rect 12102 21244 12166 21248
rect 12102 21188 12106 21244
rect 12106 21188 12162 21244
rect 12162 21188 12166 21244
rect 12102 21184 12166 21188
rect 12182 21244 12246 21248
rect 12182 21188 12186 21244
rect 12186 21188 12242 21244
rect 12242 21188 12246 21244
rect 12182 21184 12246 21188
rect 12262 21244 12326 21248
rect 12262 21188 12266 21244
rect 12266 21188 12322 21244
rect 12322 21188 12326 21244
rect 12262 21184 12326 21188
rect 23093 21244 23157 21248
rect 23093 21188 23097 21244
rect 23097 21188 23153 21244
rect 23153 21188 23157 21244
rect 23093 21184 23157 21188
rect 23173 21244 23237 21248
rect 23173 21188 23177 21244
rect 23177 21188 23233 21244
rect 23233 21188 23237 21244
rect 23173 21184 23237 21188
rect 23253 21244 23317 21248
rect 23253 21188 23257 21244
rect 23257 21188 23313 21244
rect 23313 21188 23317 21244
rect 23253 21184 23317 21188
rect 23333 21244 23397 21248
rect 23333 21188 23337 21244
rect 23337 21188 23393 21244
rect 23393 21188 23397 21244
rect 23333 21184 23397 21188
rect 6487 20700 6551 20704
rect 6487 20644 6491 20700
rect 6491 20644 6547 20700
rect 6547 20644 6551 20700
rect 6487 20640 6551 20644
rect 6567 20700 6631 20704
rect 6567 20644 6571 20700
rect 6571 20644 6627 20700
rect 6627 20644 6631 20700
rect 6567 20640 6631 20644
rect 6647 20700 6711 20704
rect 6647 20644 6651 20700
rect 6651 20644 6707 20700
rect 6707 20644 6711 20700
rect 6647 20640 6711 20644
rect 6727 20700 6791 20704
rect 6727 20644 6731 20700
rect 6731 20644 6787 20700
rect 6787 20644 6791 20700
rect 6727 20640 6791 20644
rect 17558 20700 17622 20704
rect 17558 20644 17562 20700
rect 17562 20644 17618 20700
rect 17618 20644 17622 20700
rect 17558 20640 17622 20644
rect 17638 20700 17702 20704
rect 17638 20644 17642 20700
rect 17642 20644 17698 20700
rect 17698 20644 17702 20700
rect 17638 20640 17702 20644
rect 17718 20700 17782 20704
rect 17718 20644 17722 20700
rect 17722 20644 17778 20700
rect 17778 20644 17782 20700
rect 17718 20640 17782 20644
rect 17798 20700 17862 20704
rect 17798 20644 17802 20700
rect 17802 20644 17858 20700
rect 17858 20644 17862 20700
rect 17798 20640 17862 20644
rect 28628 20700 28692 20704
rect 28628 20644 28632 20700
rect 28632 20644 28688 20700
rect 28688 20644 28692 20700
rect 28628 20640 28692 20644
rect 28708 20700 28772 20704
rect 28708 20644 28712 20700
rect 28712 20644 28768 20700
rect 28768 20644 28772 20700
rect 28708 20640 28772 20644
rect 28788 20700 28852 20704
rect 28788 20644 28792 20700
rect 28792 20644 28848 20700
rect 28848 20644 28852 20700
rect 28788 20640 28852 20644
rect 28868 20700 28932 20704
rect 28868 20644 28872 20700
rect 28872 20644 28928 20700
rect 28928 20644 28932 20700
rect 28868 20640 28932 20644
rect 12022 20156 12086 20160
rect 12022 20100 12026 20156
rect 12026 20100 12082 20156
rect 12082 20100 12086 20156
rect 12022 20096 12086 20100
rect 12102 20156 12166 20160
rect 12102 20100 12106 20156
rect 12106 20100 12162 20156
rect 12162 20100 12166 20156
rect 12102 20096 12166 20100
rect 12182 20156 12246 20160
rect 12182 20100 12186 20156
rect 12186 20100 12242 20156
rect 12242 20100 12246 20156
rect 12182 20096 12246 20100
rect 12262 20156 12326 20160
rect 12262 20100 12266 20156
rect 12266 20100 12322 20156
rect 12322 20100 12326 20156
rect 12262 20096 12326 20100
rect 23093 20156 23157 20160
rect 23093 20100 23097 20156
rect 23097 20100 23153 20156
rect 23153 20100 23157 20156
rect 23093 20096 23157 20100
rect 23173 20156 23237 20160
rect 23173 20100 23177 20156
rect 23177 20100 23233 20156
rect 23233 20100 23237 20156
rect 23173 20096 23237 20100
rect 23253 20156 23317 20160
rect 23253 20100 23257 20156
rect 23257 20100 23313 20156
rect 23313 20100 23317 20156
rect 23253 20096 23317 20100
rect 23333 20156 23397 20160
rect 23333 20100 23337 20156
rect 23337 20100 23393 20156
rect 23393 20100 23397 20156
rect 23333 20096 23397 20100
rect 6487 19612 6551 19616
rect 6487 19556 6491 19612
rect 6491 19556 6547 19612
rect 6547 19556 6551 19612
rect 6487 19552 6551 19556
rect 6567 19612 6631 19616
rect 6567 19556 6571 19612
rect 6571 19556 6627 19612
rect 6627 19556 6631 19612
rect 6567 19552 6631 19556
rect 6647 19612 6711 19616
rect 6647 19556 6651 19612
rect 6651 19556 6707 19612
rect 6707 19556 6711 19612
rect 6647 19552 6711 19556
rect 6727 19612 6791 19616
rect 6727 19556 6731 19612
rect 6731 19556 6787 19612
rect 6787 19556 6791 19612
rect 6727 19552 6791 19556
rect 17558 19612 17622 19616
rect 17558 19556 17562 19612
rect 17562 19556 17618 19612
rect 17618 19556 17622 19612
rect 17558 19552 17622 19556
rect 17638 19612 17702 19616
rect 17638 19556 17642 19612
rect 17642 19556 17698 19612
rect 17698 19556 17702 19612
rect 17638 19552 17702 19556
rect 17718 19612 17782 19616
rect 17718 19556 17722 19612
rect 17722 19556 17778 19612
rect 17778 19556 17782 19612
rect 17718 19552 17782 19556
rect 17798 19612 17862 19616
rect 17798 19556 17802 19612
rect 17802 19556 17858 19612
rect 17858 19556 17862 19612
rect 17798 19552 17862 19556
rect 28628 19612 28692 19616
rect 28628 19556 28632 19612
rect 28632 19556 28688 19612
rect 28688 19556 28692 19612
rect 28628 19552 28692 19556
rect 28708 19612 28772 19616
rect 28708 19556 28712 19612
rect 28712 19556 28768 19612
rect 28768 19556 28772 19612
rect 28708 19552 28772 19556
rect 28788 19612 28852 19616
rect 28788 19556 28792 19612
rect 28792 19556 28848 19612
rect 28848 19556 28852 19612
rect 28788 19552 28852 19556
rect 28868 19612 28932 19616
rect 28868 19556 28872 19612
rect 28872 19556 28928 19612
rect 28928 19556 28932 19612
rect 28868 19552 28932 19556
rect 12022 19068 12086 19072
rect 12022 19012 12026 19068
rect 12026 19012 12082 19068
rect 12082 19012 12086 19068
rect 12022 19008 12086 19012
rect 12102 19068 12166 19072
rect 12102 19012 12106 19068
rect 12106 19012 12162 19068
rect 12162 19012 12166 19068
rect 12102 19008 12166 19012
rect 12182 19068 12246 19072
rect 12182 19012 12186 19068
rect 12186 19012 12242 19068
rect 12242 19012 12246 19068
rect 12182 19008 12246 19012
rect 12262 19068 12326 19072
rect 12262 19012 12266 19068
rect 12266 19012 12322 19068
rect 12322 19012 12326 19068
rect 12262 19008 12326 19012
rect 23093 19068 23157 19072
rect 23093 19012 23097 19068
rect 23097 19012 23153 19068
rect 23153 19012 23157 19068
rect 23093 19008 23157 19012
rect 23173 19068 23237 19072
rect 23173 19012 23177 19068
rect 23177 19012 23233 19068
rect 23233 19012 23237 19068
rect 23173 19008 23237 19012
rect 23253 19068 23317 19072
rect 23253 19012 23257 19068
rect 23257 19012 23313 19068
rect 23313 19012 23317 19068
rect 23253 19008 23317 19012
rect 23333 19068 23397 19072
rect 23333 19012 23337 19068
rect 23337 19012 23393 19068
rect 23393 19012 23397 19068
rect 23333 19008 23397 19012
rect 6487 18524 6551 18528
rect 6487 18468 6491 18524
rect 6491 18468 6547 18524
rect 6547 18468 6551 18524
rect 6487 18464 6551 18468
rect 6567 18524 6631 18528
rect 6567 18468 6571 18524
rect 6571 18468 6627 18524
rect 6627 18468 6631 18524
rect 6567 18464 6631 18468
rect 6647 18524 6711 18528
rect 6647 18468 6651 18524
rect 6651 18468 6707 18524
rect 6707 18468 6711 18524
rect 6647 18464 6711 18468
rect 6727 18524 6791 18528
rect 6727 18468 6731 18524
rect 6731 18468 6787 18524
rect 6787 18468 6791 18524
rect 6727 18464 6791 18468
rect 17558 18524 17622 18528
rect 17558 18468 17562 18524
rect 17562 18468 17618 18524
rect 17618 18468 17622 18524
rect 17558 18464 17622 18468
rect 17638 18524 17702 18528
rect 17638 18468 17642 18524
rect 17642 18468 17698 18524
rect 17698 18468 17702 18524
rect 17638 18464 17702 18468
rect 17718 18524 17782 18528
rect 17718 18468 17722 18524
rect 17722 18468 17778 18524
rect 17778 18468 17782 18524
rect 17718 18464 17782 18468
rect 17798 18524 17862 18528
rect 17798 18468 17802 18524
rect 17802 18468 17858 18524
rect 17858 18468 17862 18524
rect 17798 18464 17862 18468
rect 28628 18524 28692 18528
rect 28628 18468 28632 18524
rect 28632 18468 28688 18524
rect 28688 18468 28692 18524
rect 28628 18464 28692 18468
rect 28708 18524 28772 18528
rect 28708 18468 28712 18524
rect 28712 18468 28768 18524
rect 28768 18468 28772 18524
rect 28708 18464 28772 18468
rect 28788 18524 28852 18528
rect 28788 18468 28792 18524
rect 28792 18468 28848 18524
rect 28848 18468 28852 18524
rect 28788 18464 28852 18468
rect 28868 18524 28932 18528
rect 28868 18468 28872 18524
rect 28872 18468 28928 18524
rect 28928 18468 28932 18524
rect 28868 18464 28932 18468
rect 12022 17980 12086 17984
rect 12022 17924 12026 17980
rect 12026 17924 12082 17980
rect 12082 17924 12086 17980
rect 12022 17920 12086 17924
rect 12102 17980 12166 17984
rect 12102 17924 12106 17980
rect 12106 17924 12162 17980
rect 12162 17924 12166 17980
rect 12102 17920 12166 17924
rect 12182 17980 12246 17984
rect 12182 17924 12186 17980
rect 12186 17924 12242 17980
rect 12242 17924 12246 17980
rect 12182 17920 12246 17924
rect 12262 17980 12326 17984
rect 12262 17924 12266 17980
rect 12266 17924 12322 17980
rect 12322 17924 12326 17980
rect 12262 17920 12326 17924
rect 23093 17980 23157 17984
rect 23093 17924 23097 17980
rect 23097 17924 23153 17980
rect 23153 17924 23157 17980
rect 23093 17920 23157 17924
rect 23173 17980 23237 17984
rect 23173 17924 23177 17980
rect 23177 17924 23233 17980
rect 23233 17924 23237 17980
rect 23173 17920 23237 17924
rect 23253 17980 23317 17984
rect 23253 17924 23257 17980
rect 23257 17924 23313 17980
rect 23313 17924 23317 17980
rect 23253 17920 23317 17924
rect 23333 17980 23397 17984
rect 23333 17924 23337 17980
rect 23337 17924 23393 17980
rect 23393 17924 23397 17980
rect 23333 17920 23397 17924
rect 6487 17436 6551 17440
rect 6487 17380 6491 17436
rect 6491 17380 6547 17436
rect 6547 17380 6551 17436
rect 6487 17376 6551 17380
rect 6567 17436 6631 17440
rect 6567 17380 6571 17436
rect 6571 17380 6627 17436
rect 6627 17380 6631 17436
rect 6567 17376 6631 17380
rect 6647 17436 6711 17440
rect 6647 17380 6651 17436
rect 6651 17380 6707 17436
rect 6707 17380 6711 17436
rect 6647 17376 6711 17380
rect 6727 17436 6791 17440
rect 6727 17380 6731 17436
rect 6731 17380 6787 17436
rect 6787 17380 6791 17436
rect 6727 17376 6791 17380
rect 17558 17436 17622 17440
rect 17558 17380 17562 17436
rect 17562 17380 17618 17436
rect 17618 17380 17622 17436
rect 17558 17376 17622 17380
rect 17638 17436 17702 17440
rect 17638 17380 17642 17436
rect 17642 17380 17698 17436
rect 17698 17380 17702 17436
rect 17638 17376 17702 17380
rect 17718 17436 17782 17440
rect 17718 17380 17722 17436
rect 17722 17380 17778 17436
rect 17778 17380 17782 17436
rect 17718 17376 17782 17380
rect 17798 17436 17862 17440
rect 17798 17380 17802 17436
rect 17802 17380 17858 17436
rect 17858 17380 17862 17436
rect 17798 17376 17862 17380
rect 28628 17436 28692 17440
rect 28628 17380 28632 17436
rect 28632 17380 28688 17436
rect 28688 17380 28692 17436
rect 28628 17376 28692 17380
rect 28708 17436 28772 17440
rect 28708 17380 28712 17436
rect 28712 17380 28768 17436
rect 28768 17380 28772 17436
rect 28708 17376 28772 17380
rect 28788 17436 28852 17440
rect 28788 17380 28792 17436
rect 28792 17380 28848 17436
rect 28848 17380 28852 17436
rect 28788 17376 28852 17380
rect 28868 17436 28932 17440
rect 28868 17380 28872 17436
rect 28872 17380 28928 17436
rect 28928 17380 28932 17436
rect 28868 17376 28932 17380
rect 12022 16892 12086 16896
rect 12022 16836 12026 16892
rect 12026 16836 12082 16892
rect 12082 16836 12086 16892
rect 12022 16832 12086 16836
rect 12102 16892 12166 16896
rect 12102 16836 12106 16892
rect 12106 16836 12162 16892
rect 12162 16836 12166 16892
rect 12102 16832 12166 16836
rect 12182 16892 12246 16896
rect 12182 16836 12186 16892
rect 12186 16836 12242 16892
rect 12242 16836 12246 16892
rect 12182 16832 12246 16836
rect 12262 16892 12326 16896
rect 12262 16836 12266 16892
rect 12266 16836 12322 16892
rect 12322 16836 12326 16892
rect 12262 16832 12326 16836
rect 23093 16892 23157 16896
rect 23093 16836 23097 16892
rect 23097 16836 23153 16892
rect 23153 16836 23157 16892
rect 23093 16832 23157 16836
rect 23173 16892 23237 16896
rect 23173 16836 23177 16892
rect 23177 16836 23233 16892
rect 23233 16836 23237 16892
rect 23173 16832 23237 16836
rect 23253 16892 23317 16896
rect 23253 16836 23257 16892
rect 23257 16836 23313 16892
rect 23313 16836 23317 16892
rect 23253 16832 23317 16836
rect 23333 16892 23397 16896
rect 23333 16836 23337 16892
rect 23337 16836 23393 16892
rect 23393 16836 23397 16892
rect 23333 16832 23397 16836
rect 6487 16348 6551 16352
rect 6487 16292 6491 16348
rect 6491 16292 6547 16348
rect 6547 16292 6551 16348
rect 6487 16288 6551 16292
rect 6567 16348 6631 16352
rect 6567 16292 6571 16348
rect 6571 16292 6627 16348
rect 6627 16292 6631 16348
rect 6567 16288 6631 16292
rect 6647 16348 6711 16352
rect 6647 16292 6651 16348
rect 6651 16292 6707 16348
rect 6707 16292 6711 16348
rect 6647 16288 6711 16292
rect 6727 16348 6791 16352
rect 6727 16292 6731 16348
rect 6731 16292 6787 16348
rect 6787 16292 6791 16348
rect 6727 16288 6791 16292
rect 17558 16348 17622 16352
rect 17558 16292 17562 16348
rect 17562 16292 17618 16348
rect 17618 16292 17622 16348
rect 17558 16288 17622 16292
rect 17638 16348 17702 16352
rect 17638 16292 17642 16348
rect 17642 16292 17698 16348
rect 17698 16292 17702 16348
rect 17638 16288 17702 16292
rect 17718 16348 17782 16352
rect 17718 16292 17722 16348
rect 17722 16292 17778 16348
rect 17778 16292 17782 16348
rect 17718 16288 17782 16292
rect 17798 16348 17862 16352
rect 17798 16292 17802 16348
rect 17802 16292 17858 16348
rect 17858 16292 17862 16348
rect 17798 16288 17862 16292
rect 28628 16348 28692 16352
rect 28628 16292 28632 16348
rect 28632 16292 28688 16348
rect 28688 16292 28692 16348
rect 28628 16288 28692 16292
rect 28708 16348 28772 16352
rect 28708 16292 28712 16348
rect 28712 16292 28768 16348
rect 28768 16292 28772 16348
rect 28708 16288 28772 16292
rect 28788 16348 28852 16352
rect 28788 16292 28792 16348
rect 28792 16292 28848 16348
rect 28848 16292 28852 16348
rect 28788 16288 28852 16292
rect 28868 16348 28932 16352
rect 28868 16292 28872 16348
rect 28872 16292 28928 16348
rect 28928 16292 28932 16348
rect 28868 16288 28932 16292
rect 12022 15804 12086 15808
rect 12022 15748 12026 15804
rect 12026 15748 12082 15804
rect 12082 15748 12086 15804
rect 12022 15744 12086 15748
rect 12102 15804 12166 15808
rect 12102 15748 12106 15804
rect 12106 15748 12162 15804
rect 12162 15748 12166 15804
rect 12102 15744 12166 15748
rect 12182 15804 12246 15808
rect 12182 15748 12186 15804
rect 12186 15748 12242 15804
rect 12242 15748 12246 15804
rect 12182 15744 12246 15748
rect 12262 15804 12326 15808
rect 12262 15748 12266 15804
rect 12266 15748 12322 15804
rect 12322 15748 12326 15804
rect 12262 15744 12326 15748
rect 23093 15804 23157 15808
rect 23093 15748 23097 15804
rect 23097 15748 23153 15804
rect 23153 15748 23157 15804
rect 23093 15744 23157 15748
rect 23173 15804 23237 15808
rect 23173 15748 23177 15804
rect 23177 15748 23233 15804
rect 23233 15748 23237 15804
rect 23173 15744 23237 15748
rect 23253 15804 23317 15808
rect 23253 15748 23257 15804
rect 23257 15748 23313 15804
rect 23313 15748 23317 15804
rect 23253 15744 23317 15748
rect 23333 15804 23397 15808
rect 23333 15748 23337 15804
rect 23337 15748 23393 15804
rect 23393 15748 23397 15804
rect 23333 15744 23397 15748
rect 6487 15260 6551 15264
rect 6487 15204 6491 15260
rect 6491 15204 6547 15260
rect 6547 15204 6551 15260
rect 6487 15200 6551 15204
rect 6567 15260 6631 15264
rect 6567 15204 6571 15260
rect 6571 15204 6627 15260
rect 6627 15204 6631 15260
rect 6567 15200 6631 15204
rect 6647 15260 6711 15264
rect 6647 15204 6651 15260
rect 6651 15204 6707 15260
rect 6707 15204 6711 15260
rect 6647 15200 6711 15204
rect 6727 15260 6791 15264
rect 6727 15204 6731 15260
rect 6731 15204 6787 15260
rect 6787 15204 6791 15260
rect 6727 15200 6791 15204
rect 17558 15260 17622 15264
rect 17558 15204 17562 15260
rect 17562 15204 17618 15260
rect 17618 15204 17622 15260
rect 17558 15200 17622 15204
rect 17638 15260 17702 15264
rect 17638 15204 17642 15260
rect 17642 15204 17698 15260
rect 17698 15204 17702 15260
rect 17638 15200 17702 15204
rect 17718 15260 17782 15264
rect 17718 15204 17722 15260
rect 17722 15204 17778 15260
rect 17778 15204 17782 15260
rect 17718 15200 17782 15204
rect 17798 15260 17862 15264
rect 17798 15204 17802 15260
rect 17802 15204 17858 15260
rect 17858 15204 17862 15260
rect 17798 15200 17862 15204
rect 28628 15260 28692 15264
rect 28628 15204 28632 15260
rect 28632 15204 28688 15260
rect 28688 15204 28692 15260
rect 28628 15200 28692 15204
rect 28708 15260 28772 15264
rect 28708 15204 28712 15260
rect 28712 15204 28768 15260
rect 28768 15204 28772 15260
rect 28708 15200 28772 15204
rect 28788 15260 28852 15264
rect 28788 15204 28792 15260
rect 28792 15204 28848 15260
rect 28848 15204 28852 15260
rect 28788 15200 28852 15204
rect 28868 15260 28932 15264
rect 28868 15204 28872 15260
rect 28872 15204 28928 15260
rect 28928 15204 28932 15260
rect 28868 15200 28932 15204
rect 12022 14716 12086 14720
rect 12022 14660 12026 14716
rect 12026 14660 12082 14716
rect 12082 14660 12086 14716
rect 12022 14656 12086 14660
rect 12102 14716 12166 14720
rect 12102 14660 12106 14716
rect 12106 14660 12162 14716
rect 12162 14660 12166 14716
rect 12102 14656 12166 14660
rect 12182 14716 12246 14720
rect 12182 14660 12186 14716
rect 12186 14660 12242 14716
rect 12242 14660 12246 14716
rect 12182 14656 12246 14660
rect 12262 14716 12326 14720
rect 12262 14660 12266 14716
rect 12266 14660 12322 14716
rect 12322 14660 12326 14716
rect 12262 14656 12326 14660
rect 23093 14716 23157 14720
rect 23093 14660 23097 14716
rect 23097 14660 23153 14716
rect 23153 14660 23157 14716
rect 23093 14656 23157 14660
rect 23173 14716 23237 14720
rect 23173 14660 23177 14716
rect 23177 14660 23233 14716
rect 23233 14660 23237 14716
rect 23173 14656 23237 14660
rect 23253 14716 23317 14720
rect 23253 14660 23257 14716
rect 23257 14660 23313 14716
rect 23313 14660 23317 14716
rect 23253 14656 23317 14660
rect 23333 14716 23397 14720
rect 23333 14660 23337 14716
rect 23337 14660 23393 14716
rect 23393 14660 23397 14716
rect 23333 14656 23397 14660
rect 6487 14172 6551 14176
rect 6487 14116 6491 14172
rect 6491 14116 6547 14172
rect 6547 14116 6551 14172
rect 6487 14112 6551 14116
rect 6567 14172 6631 14176
rect 6567 14116 6571 14172
rect 6571 14116 6627 14172
rect 6627 14116 6631 14172
rect 6567 14112 6631 14116
rect 6647 14172 6711 14176
rect 6647 14116 6651 14172
rect 6651 14116 6707 14172
rect 6707 14116 6711 14172
rect 6647 14112 6711 14116
rect 6727 14172 6791 14176
rect 6727 14116 6731 14172
rect 6731 14116 6787 14172
rect 6787 14116 6791 14172
rect 6727 14112 6791 14116
rect 17558 14172 17622 14176
rect 17558 14116 17562 14172
rect 17562 14116 17618 14172
rect 17618 14116 17622 14172
rect 17558 14112 17622 14116
rect 17638 14172 17702 14176
rect 17638 14116 17642 14172
rect 17642 14116 17698 14172
rect 17698 14116 17702 14172
rect 17638 14112 17702 14116
rect 17718 14172 17782 14176
rect 17718 14116 17722 14172
rect 17722 14116 17778 14172
rect 17778 14116 17782 14172
rect 17718 14112 17782 14116
rect 17798 14172 17862 14176
rect 17798 14116 17802 14172
rect 17802 14116 17858 14172
rect 17858 14116 17862 14172
rect 17798 14112 17862 14116
rect 28628 14172 28692 14176
rect 28628 14116 28632 14172
rect 28632 14116 28688 14172
rect 28688 14116 28692 14172
rect 28628 14112 28692 14116
rect 28708 14172 28772 14176
rect 28708 14116 28712 14172
rect 28712 14116 28768 14172
rect 28768 14116 28772 14172
rect 28708 14112 28772 14116
rect 28788 14172 28852 14176
rect 28788 14116 28792 14172
rect 28792 14116 28848 14172
rect 28848 14116 28852 14172
rect 28788 14112 28852 14116
rect 28868 14172 28932 14176
rect 28868 14116 28872 14172
rect 28872 14116 28928 14172
rect 28928 14116 28932 14172
rect 28868 14112 28932 14116
rect 12022 13628 12086 13632
rect 12022 13572 12026 13628
rect 12026 13572 12082 13628
rect 12082 13572 12086 13628
rect 12022 13568 12086 13572
rect 12102 13628 12166 13632
rect 12102 13572 12106 13628
rect 12106 13572 12162 13628
rect 12162 13572 12166 13628
rect 12102 13568 12166 13572
rect 12182 13628 12246 13632
rect 12182 13572 12186 13628
rect 12186 13572 12242 13628
rect 12242 13572 12246 13628
rect 12182 13568 12246 13572
rect 12262 13628 12326 13632
rect 12262 13572 12266 13628
rect 12266 13572 12322 13628
rect 12322 13572 12326 13628
rect 12262 13568 12326 13572
rect 23093 13628 23157 13632
rect 23093 13572 23097 13628
rect 23097 13572 23153 13628
rect 23153 13572 23157 13628
rect 23093 13568 23157 13572
rect 23173 13628 23237 13632
rect 23173 13572 23177 13628
rect 23177 13572 23233 13628
rect 23233 13572 23237 13628
rect 23173 13568 23237 13572
rect 23253 13628 23317 13632
rect 23253 13572 23257 13628
rect 23257 13572 23313 13628
rect 23313 13572 23317 13628
rect 23253 13568 23317 13572
rect 23333 13628 23397 13632
rect 23333 13572 23337 13628
rect 23337 13572 23393 13628
rect 23393 13572 23397 13628
rect 23333 13568 23397 13572
rect 6487 13084 6551 13088
rect 6487 13028 6491 13084
rect 6491 13028 6547 13084
rect 6547 13028 6551 13084
rect 6487 13024 6551 13028
rect 6567 13084 6631 13088
rect 6567 13028 6571 13084
rect 6571 13028 6627 13084
rect 6627 13028 6631 13084
rect 6567 13024 6631 13028
rect 6647 13084 6711 13088
rect 6647 13028 6651 13084
rect 6651 13028 6707 13084
rect 6707 13028 6711 13084
rect 6647 13024 6711 13028
rect 6727 13084 6791 13088
rect 6727 13028 6731 13084
rect 6731 13028 6787 13084
rect 6787 13028 6791 13084
rect 6727 13024 6791 13028
rect 17558 13084 17622 13088
rect 17558 13028 17562 13084
rect 17562 13028 17618 13084
rect 17618 13028 17622 13084
rect 17558 13024 17622 13028
rect 17638 13084 17702 13088
rect 17638 13028 17642 13084
rect 17642 13028 17698 13084
rect 17698 13028 17702 13084
rect 17638 13024 17702 13028
rect 17718 13084 17782 13088
rect 17718 13028 17722 13084
rect 17722 13028 17778 13084
rect 17778 13028 17782 13084
rect 17718 13024 17782 13028
rect 17798 13084 17862 13088
rect 17798 13028 17802 13084
rect 17802 13028 17858 13084
rect 17858 13028 17862 13084
rect 17798 13024 17862 13028
rect 28628 13084 28692 13088
rect 28628 13028 28632 13084
rect 28632 13028 28688 13084
rect 28688 13028 28692 13084
rect 28628 13024 28692 13028
rect 28708 13084 28772 13088
rect 28708 13028 28712 13084
rect 28712 13028 28768 13084
rect 28768 13028 28772 13084
rect 28708 13024 28772 13028
rect 28788 13084 28852 13088
rect 28788 13028 28792 13084
rect 28792 13028 28848 13084
rect 28848 13028 28852 13084
rect 28788 13024 28852 13028
rect 28868 13084 28932 13088
rect 28868 13028 28872 13084
rect 28872 13028 28928 13084
rect 28928 13028 28932 13084
rect 28868 13024 28932 13028
rect 12022 12540 12086 12544
rect 12022 12484 12026 12540
rect 12026 12484 12082 12540
rect 12082 12484 12086 12540
rect 12022 12480 12086 12484
rect 12102 12540 12166 12544
rect 12102 12484 12106 12540
rect 12106 12484 12162 12540
rect 12162 12484 12166 12540
rect 12102 12480 12166 12484
rect 12182 12540 12246 12544
rect 12182 12484 12186 12540
rect 12186 12484 12242 12540
rect 12242 12484 12246 12540
rect 12182 12480 12246 12484
rect 12262 12540 12326 12544
rect 12262 12484 12266 12540
rect 12266 12484 12322 12540
rect 12322 12484 12326 12540
rect 12262 12480 12326 12484
rect 23093 12540 23157 12544
rect 23093 12484 23097 12540
rect 23097 12484 23153 12540
rect 23153 12484 23157 12540
rect 23093 12480 23157 12484
rect 23173 12540 23237 12544
rect 23173 12484 23177 12540
rect 23177 12484 23233 12540
rect 23233 12484 23237 12540
rect 23173 12480 23237 12484
rect 23253 12540 23317 12544
rect 23253 12484 23257 12540
rect 23257 12484 23313 12540
rect 23313 12484 23317 12540
rect 23253 12480 23317 12484
rect 23333 12540 23397 12544
rect 23333 12484 23337 12540
rect 23337 12484 23393 12540
rect 23393 12484 23397 12540
rect 23333 12480 23397 12484
rect 6487 11996 6551 12000
rect 6487 11940 6491 11996
rect 6491 11940 6547 11996
rect 6547 11940 6551 11996
rect 6487 11936 6551 11940
rect 6567 11996 6631 12000
rect 6567 11940 6571 11996
rect 6571 11940 6627 11996
rect 6627 11940 6631 11996
rect 6567 11936 6631 11940
rect 6647 11996 6711 12000
rect 6647 11940 6651 11996
rect 6651 11940 6707 11996
rect 6707 11940 6711 11996
rect 6647 11936 6711 11940
rect 6727 11996 6791 12000
rect 6727 11940 6731 11996
rect 6731 11940 6787 11996
rect 6787 11940 6791 11996
rect 6727 11936 6791 11940
rect 17558 11996 17622 12000
rect 17558 11940 17562 11996
rect 17562 11940 17618 11996
rect 17618 11940 17622 11996
rect 17558 11936 17622 11940
rect 17638 11996 17702 12000
rect 17638 11940 17642 11996
rect 17642 11940 17698 11996
rect 17698 11940 17702 11996
rect 17638 11936 17702 11940
rect 17718 11996 17782 12000
rect 17718 11940 17722 11996
rect 17722 11940 17778 11996
rect 17778 11940 17782 11996
rect 17718 11936 17782 11940
rect 17798 11996 17862 12000
rect 17798 11940 17802 11996
rect 17802 11940 17858 11996
rect 17858 11940 17862 11996
rect 17798 11936 17862 11940
rect 28628 11996 28692 12000
rect 28628 11940 28632 11996
rect 28632 11940 28688 11996
rect 28688 11940 28692 11996
rect 28628 11936 28692 11940
rect 28708 11996 28772 12000
rect 28708 11940 28712 11996
rect 28712 11940 28768 11996
rect 28768 11940 28772 11996
rect 28708 11936 28772 11940
rect 28788 11996 28852 12000
rect 28788 11940 28792 11996
rect 28792 11940 28848 11996
rect 28848 11940 28852 11996
rect 28788 11936 28852 11940
rect 28868 11996 28932 12000
rect 28868 11940 28872 11996
rect 28872 11940 28928 11996
rect 28928 11940 28932 11996
rect 28868 11936 28932 11940
rect 12022 11452 12086 11456
rect 12022 11396 12026 11452
rect 12026 11396 12082 11452
rect 12082 11396 12086 11452
rect 12022 11392 12086 11396
rect 12102 11452 12166 11456
rect 12102 11396 12106 11452
rect 12106 11396 12162 11452
rect 12162 11396 12166 11452
rect 12102 11392 12166 11396
rect 12182 11452 12246 11456
rect 12182 11396 12186 11452
rect 12186 11396 12242 11452
rect 12242 11396 12246 11452
rect 12182 11392 12246 11396
rect 12262 11452 12326 11456
rect 12262 11396 12266 11452
rect 12266 11396 12322 11452
rect 12322 11396 12326 11452
rect 12262 11392 12326 11396
rect 23093 11452 23157 11456
rect 23093 11396 23097 11452
rect 23097 11396 23153 11452
rect 23153 11396 23157 11452
rect 23093 11392 23157 11396
rect 23173 11452 23237 11456
rect 23173 11396 23177 11452
rect 23177 11396 23233 11452
rect 23233 11396 23237 11452
rect 23173 11392 23237 11396
rect 23253 11452 23317 11456
rect 23253 11396 23257 11452
rect 23257 11396 23313 11452
rect 23313 11396 23317 11452
rect 23253 11392 23317 11396
rect 23333 11452 23397 11456
rect 23333 11396 23337 11452
rect 23337 11396 23393 11452
rect 23393 11396 23397 11452
rect 23333 11392 23397 11396
rect 6487 10908 6551 10912
rect 6487 10852 6491 10908
rect 6491 10852 6547 10908
rect 6547 10852 6551 10908
rect 6487 10848 6551 10852
rect 6567 10908 6631 10912
rect 6567 10852 6571 10908
rect 6571 10852 6627 10908
rect 6627 10852 6631 10908
rect 6567 10848 6631 10852
rect 6647 10908 6711 10912
rect 6647 10852 6651 10908
rect 6651 10852 6707 10908
rect 6707 10852 6711 10908
rect 6647 10848 6711 10852
rect 6727 10908 6791 10912
rect 6727 10852 6731 10908
rect 6731 10852 6787 10908
rect 6787 10852 6791 10908
rect 6727 10848 6791 10852
rect 17558 10908 17622 10912
rect 17558 10852 17562 10908
rect 17562 10852 17618 10908
rect 17618 10852 17622 10908
rect 17558 10848 17622 10852
rect 17638 10908 17702 10912
rect 17638 10852 17642 10908
rect 17642 10852 17698 10908
rect 17698 10852 17702 10908
rect 17638 10848 17702 10852
rect 17718 10908 17782 10912
rect 17718 10852 17722 10908
rect 17722 10852 17778 10908
rect 17778 10852 17782 10908
rect 17718 10848 17782 10852
rect 17798 10908 17862 10912
rect 17798 10852 17802 10908
rect 17802 10852 17858 10908
rect 17858 10852 17862 10908
rect 17798 10848 17862 10852
rect 28628 10908 28692 10912
rect 28628 10852 28632 10908
rect 28632 10852 28688 10908
rect 28688 10852 28692 10908
rect 28628 10848 28692 10852
rect 28708 10908 28772 10912
rect 28708 10852 28712 10908
rect 28712 10852 28768 10908
rect 28768 10852 28772 10908
rect 28708 10848 28772 10852
rect 28788 10908 28852 10912
rect 28788 10852 28792 10908
rect 28792 10852 28848 10908
rect 28848 10852 28852 10908
rect 28788 10848 28852 10852
rect 28868 10908 28932 10912
rect 28868 10852 28872 10908
rect 28872 10852 28928 10908
rect 28928 10852 28932 10908
rect 28868 10848 28932 10852
rect 12022 10364 12086 10368
rect 12022 10308 12026 10364
rect 12026 10308 12082 10364
rect 12082 10308 12086 10364
rect 12022 10304 12086 10308
rect 12102 10364 12166 10368
rect 12102 10308 12106 10364
rect 12106 10308 12162 10364
rect 12162 10308 12166 10364
rect 12102 10304 12166 10308
rect 12182 10364 12246 10368
rect 12182 10308 12186 10364
rect 12186 10308 12242 10364
rect 12242 10308 12246 10364
rect 12182 10304 12246 10308
rect 12262 10364 12326 10368
rect 12262 10308 12266 10364
rect 12266 10308 12322 10364
rect 12322 10308 12326 10364
rect 12262 10304 12326 10308
rect 23093 10364 23157 10368
rect 23093 10308 23097 10364
rect 23097 10308 23153 10364
rect 23153 10308 23157 10364
rect 23093 10304 23157 10308
rect 23173 10364 23237 10368
rect 23173 10308 23177 10364
rect 23177 10308 23233 10364
rect 23233 10308 23237 10364
rect 23173 10304 23237 10308
rect 23253 10364 23317 10368
rect 23253 10308 23257 10364
rect 23257 10308 23313 10364
rect 23313 10308 23317 10364
rect 23253 10304 23317 10308
rect 23333 10364 23397 10368
rect 23333 10308 23337 10364
rect 23337 10308 23393 10364
rect 23393 10308 23397 10364
rect 23333 10304 23397 10308
rect 6487 9820 6551 9824
rect 6487 9764 6491 9820
rect 6491 9764 6547 9820
rect 6547 9764 6551 9820
rect 6487 9760 6551 9764
rect 6567 9820 6631 9824
rect 6567 9764 6571 9820
rect 6571 9764 6627 9820
rect 6627 9764 6631 9820
rect 6567 9760 6631 9764
rect 6647 9820 6711 9824
rect 6647 9764 6651 9820
rect 6651 9764 6707 9820
rect 6707 9764 6711 9820
rect 6647 9760 6711 9764
rect 6727 9820 6791 9824
rect 6727 9764 6731 9820
rect 6731 9764 6787 9820
rect 6787 9764 6791 9820
rect 6727 9760 6791 9764
rect 17558 9820 17622 9824
rect 17558 9764 17562 9820
rect 17562 9764 17618 9820
rect 17618 9764 17622 9820
rect 17558 9760 17622 9764
rect 17638 9820 17702 9824
rect 17638 9764 17642 9820
rect 17642 9764 17698 9820
rect 17698 9764 17702 9820
rect 17638 9760 17702 9764
rect 17718 9820 17782 9824
rect 17718 9764 17722 9820
rect 17722 9764 17778 9820
rect 17778 9764 17782 9820
rect 17718 9760 17782 9764
rect 17798 9820 17862 9824
rect 17798 9764 17802 9820
rect 17802 9764 17858 9820
rect 17858 9764 17862 9820
rect 17798 9760 17862 9764
rect 28628 9820 28692 9824
rect 28628 9764 28632 9820
rect 28632 9764 28688 9820
rect 28688 9764 28692 9820
rect 28628 9760 28692 9764
rect 28708 9820 28772 9824
rect 28708 9764 28712 9820
rect 28712 9764 28768 9820
rect 28768 9764 28772 9820
rect 28708 9760 28772 9764
rect 28788 9820 28852 9824
rect 28788 9764 28792 9820
rect 28792 9764 28848 9820
rect 28848 9764 28852 9820
rect 28788 9760 28852 9764
rect 28868 9820 28932 9824
rect 28868 9764 28872 9820
rect 28872 9764 28928 9820
rect 28928 9764 28932 9820
rect 28868 9760 28932 9764
rect 12022 9276 12086 9280
rect 12022 9220 12026 9276
rect 12026 9220 12082 9276
rect 12082 9220 12086 9276
rect 12022 9216 12086 9220
rect 12102 9276 12166 9280
rect 12102 9220 12106 9276
rect 12106 9220 12162 9276
rect 12162 9220 12166 9276
rect 12102 9216 12166 9220
rect 12182 9276 12246 9280
rect 12182 9220 12186 9276
rect 12186 9220 12242 9276
rect 12242 9220 12246 9276
rect 12182 9216 12246 9220
rect 12262 9276 12326 9280
rect 12262 9220 12266 9276
rect 12266 9220 12322 9276
rect 12322 9220 12326 9276
rect 12262 9216 12326 9220
rect 23093 9276 23157 9280
rect 23093 9220 23097 9276
rect 23097 9220 23153 9276
rect 23153 9220 23157 9276
rect 23093 9216 23157 9220
rect 23173 9276 23237 9280
rect 23173 9220 23177 9276
rect 23177 9220 23233 9276
rect 23233 9220 23237 9276
rect 23173 9216 23237 9220
rect 23253 9276 23317 9280
rect 23253 9220 23257 9276
rect 23257 9220 23313 9276
rect 23313 9220 23317 9276
rect 23253 9216 23317 9220
rect 23333 9276 23397 9280
rect 23333 9220 23337 9276
rect 23337 9220 23393 9276
rect 23393 9220 23397 9276
rect 23333 9216 23397 9220
rect 6487 8732 6551 8736
rect 6487 8676 6491 8732
rect 6491 8676 6547 8732
rect 6547 8676 6551 8732
rect 6487 8672 6551 8676
rect 6567 8732 6631 8736
rect 6567 8676 6571 8732
rect 6571 8676 6627 8732
rect 6627 8676 6631 8732
rect 6567 8672 6631 8676
rect 6647 8732 6711 8736
rect 6647 8676 6651 8732
rect 6651 8676 6707 8732
rect 6707 8676 6711 8732
rect 6647 8672 6711 8676
rect 6727 8732 6791 8736
rect 6727 8676 6731 8732
rect 6731 8676 6787 8732
rect 6787 8676 6791 8732
rect 6727 8672 6791 8676
rect 17558 8732 17622 8736
rect 17558 8676 17562 8732
rect 17562 8676 17618 8732
rect 17618 8676 17622 8732
rect 17558 8672 17622 8676
rect 17638 8732 17702 8736
rect 17638 8676 17642 8732
rect 17642 8676 17698 8732
rect 17698 8676 17702 8732
rect 17638 8672 17702 8676
rect 17718 8732 17782 8736
rect 17718 8676 17722 8732
rect 17722 8676 17778 8732
rect 17778 8676 17782 8732
rect 17718 8672 17782 8676
rect 17798 8732 17862 8736
rect 17798 8676 17802 8732
rect 17802 8676 17858 8732
rect 17858 8676 17862 8732
rect 17798 8672 17862 8676
rect 28628 8732 28692 8736
rect 28628 8676 28632 8732
rect 28632 8676 28688 8732
rect 28688 8676 28692 8732
rect 28628 8672 28692 8676
rect 28708 8732 28772 8736
rect 28708 8676 28712 8732
rect 28712 8676 28768 8732
rect 28768 8676 28772 8732
rect 28708 8672 28772 8676
rect 28788 8732 28852 8736
rect 28788 8676 28792 8732
rect 28792 8676 28848 8732
rect 28848 8676 28852 8732
rect 28788 8672 28852 8676
rect 28868 8732 28932 8736
rect 28868 8676 28872 8732
rect 28872 8676 28928 8732
rect 28928 8676 28932 8732
rect 28868 8672 28932 8676
rect 12022 8188 12086 8192
rect 12022 8132 12026 8188
rect 12026 8132 12082 8188
rect 12082 8132 12086 8188
rect 12022 8128 12086 8132
rect 12102 8188 12166 8192
rect 12102 8132 12106 8188
rect 12106 8132 12162 8188
rect 12162 8132 12166 8188
rect 12102 8128 12166 8132
rect 12182 8188 12246 8192
rect 12182 8132 12186 8188
rect 12186 8132 12242 8188
rect 12242 8132 12246 8188
rect 12182 8128 12246 8132
rect 12262 8188 12326 8192
rect 12262 8132 12266 8188
rect 12266 8132 12322 8188
rect 12322 8132 12326 8188
rect 12262 8128 12326 8132
rect 23093 8188 23157 8192
rect 23093 8132 23097 8188
rect 23097 8132 23153 8188
rect 23153 8132 23157 8188
rect 23093 8128 23157 8132
rect 23173 8188 23237 8192
rect 23173 8132 23177 8188
rect 23177 8132 23233 8188
rect 23233 8132 23237 8188
rect 23173 8128 23237 8132
rect 23253 8188 23317 8192
rect 23253 8132 23257 8188
rect 23257 8132 23313 8188
rect 23313 8132 23317 8188
rect 23253 8128 23317 8132
rect 23333 8188 23397 8192
rect 23333 8132 23337 8188
rect 23337 8132 23393 8188
rect 23393 8132 23397 8188
rect 23333 8128 23397 8132
rect 6487 7644 6551 7648
rect 6487 7588 6491 7644
rect 6491 7588 6547 7644
rect 6547 7588 6551 7644
rect 6487 7584 6551 7588
rect 6567 7644 6631 7648
rect 6567 7588 6571 7644
rect 6571 7588 6627 7644
rect 6627 7588 6631 7644
rect 6567 7584 6631 7588
rect 6647 7644 6711 7648
rect 6647 7588 6651 7644
rect 6651 7588 6707 7644
rect 6707 7588 6711 7644
rect 6647 7584 6711 7588
rect 6727 7644 6791 7648
rect 6727 7588 6731 7644
rect 6731 7588 6787 7644
rect 6787 7588 6791 7644
rect 6727 7584 6791 7588
rect 17558 7644 17622 7648
rect 17558 7588 17562 7644
rect 17562 7588 17618 7644
rect 17618 7588 17622 7644
rect 17558 7584 17622 7588
rect 17638 7644 17702 7648
rect 17638 7588 17642 7644
rect 17642 7588 17698 7644
rect 17698 7588 17702 7644
rect 17638 7584 17702 7588
rect 17718 7644 17782 7648
rect 17718 7588 17722 7644
rect 17722 7588 17778 7644
rect 17778 7588 17782 7644
rect 17718 7584 17782 7588
rect 17798 7644 17862 7648
rect 17798 7588 17802 7644
rect 17802 7588 17858 7644
rect 17858 7588 17862 7644
rect 17798 7584 17862 7588
rect 28628 7644 28692 7648
rect 28628 7588 28632 7644
rect 28632 7588 28688 7644
rect 28688 7588 28692 7644
rect 28628 7584 28692 7588
rect 28708 7644 28772 7648
rect 28708 7588 28712 7644
rect 28712 7588 28768 7644
rect 28768 7588 28772 7644
rect 28708 7584 28772 7588
rect 28788 7644 28852 7648
rect 28788 7588 28792 7644
rect 28792 7588 28848 7644
rect 28848 7588 28852 7644
rect 28788 7584 28852 7588
rect 28868 7644 28932 7648
rect 28868 7588 28872 7644
rect 28872 7588 28928 7644
rect 28928 7588 28932 7644
rect 28868 7584 28932 7588
rect 12022 7100 12086 7104
rect 12022 7044 12026 7100
rect 12026 7044 12082 7100
rect 12082 7044 12086 7100
rect 12022 7040 12086 7044
rect 12102 7100 12166 7104
rect 12102 7044 12106 7100
rect 12106 7044 12162 7100
rect 12162 7044 12166 7100
rect 12102 7040 12166 7044
rect 12182 7100 12246 7104
rect 12182 7044 12186 7100
rect 12186 7044 12242 7100
rect 12242 7044 12246 7100
rect 12182 7040 12246 7044
rect 12262 7100 12326 7104
rect 12262 7044 12266 7100
rect 12266 7044 12322 7100
rect 12322 7044 12326 7100
rect 12262 7040 12326 7044
rect 23093 7100 23157 7104
rect 23093 7044 23097 7100
rect 23097 7044 23153 7100
rect 23153 7044 23157 7100
rect 23093 7040 23157 7044
rect 23173 7100 23237 7104
rect 23173 7044 23177 7100
rect 23177 7044 23233 7100
rect 23233 7044 23237 7100
rect 23173 7040 23237 7044
rect 23253 7100 23317 7104
rect 23253 7044 23257 7100
rect 23257 7044 23313 7100
rect 23313 7044 23317 7100
rect 23253 7040 23317 7044
rect 23333 7100 23397 7104
rect 23333 7044 23337 7100
rect 23337 7044 23393 7100
rect 23393 7044 23397 7100
rect 23333 7040 23397 7044
rect 6487 6556 6551 6560
rect 6487 6500 6491 6556
rect 6491 6500 6547 6556
rect 6547 6500 6551 6556
rect 6487 6496 6551 6500
rect 6567 6556 6631 6560
rect 6567 6500 6571 6556
rect 6571 6500 6627 6556
rect 6627 6500 6631 6556
rect 6567 6496 6631 6500
rect 6647 6556 6711 6560
rect 6647 6500 6651 6556
rect 6651 6500 6707 6556
rect 6707 6500 6711 6556
rect 6647 6496 6711 6500
rect 6727 6556 6791 6560
rect 6727 6500 6731 6556
rect 6731 6500 6787 6556
rect 6787 6500 6791 6556
rect 6727 6496 6791 6500
rect 17558 6556 17622 6560
rect 17558 6500 17562 6556
rect 17562 6500 17618 6556
rect 17618 6500 17622 6556
rect 17558 6496 17622 6500
rect 17638 6556 17702 6560
rect 17638 6500 17642 6556
rect 17642 6500 17698 6556
rect 17698 6500 17702 6556
rect 17638 6496 17702 6500
rect 17718 6556 17782 6560
rect 17718 6500 17722 6556
rect 17722 6500 17778 6556
rect 17778 6500 17782 6556
rect 17718 6496 17782 6500
rect 17798 6556 17862 6560
rect 17798 6500 17802 6556
rect 17802 6500 17858 6556
rect 17858 6500 17862 6556
rect 17798 6496 17862 6500
rect 28628 6556 28692 6560
rect 28628 6500 28632 6556
rect 28632 6500 28688 6556
rect 28688 6500 28692 6556
rect 28628 6496 28692 6500
rect 28708 6556 28772 6560
rect 28708 6500 28712 6556
rect 28712 6500 28768 6556
rect 28768 6500 28772 6556
rect 28708 6496 28772 6500
rect 28788 6556 28852 6560
rect 28788 6500 28792 6556
rect 28792 6500 28848 6556
rect 28848 6500 28852 6556
rect 28788 6496 28852 6500
rect 28868 6556 28932 6560
rect 28868 6500 28872 6556
rect 28872 6500 28928 6556
rect 28928 6500 28932 6556
rect 28868 6496 28932 6500
rect 12022 6012 12086 6016
rect 12022 5956 12026 6012
rect 12026 5956 12082 6012
rect 12082 5956 12086 6012
rect 12022 5952 12086 5956
rect 12102 6012 12166 6016
rect 12102 5956 12106 6012
rect 12106 5956 12162 6012
rect 12162 5956 12166 6012
rect 12102 5952 12166 5956
rect 12182 6012 12246 6016
rect 12182 5956 12186 6012
rect 12186 5956 12242 6012
rect 12242 5956 12246 6012
rect 12182 5952 12246 5956
rect 12262 6012 12326 6016
rect 12262 5956 12266 6012
rect 12266 5956 12322 6012
rect 12322 5956 12326 6012
rect 12262 5952 12326 5956
rect 23093 6012 23157 6016
rect 23093 5956 23097 6012
rect 23097 5956 23153 6012
rect 23153 5956 23157 6012
rect 23093 5952 23157 5956
rect 23173 6012 23237 6016
rect 23173 5956 23177 6012
rect 23177 5956 23233 6012
rect 23233 5956 23237 6012
rect 23173 5952 23237 5956
rect 23253 6012 23317 6016
rect 23253 5956 23257 6012
rect 23257 5956 23313 6012
rect 23313 5956 23317 6012
rect 23253 5952 23317 5956
rect 23333 6012 23397 6016
rect 23333 5956 23337 6012
rect 23337 5956 23393 6012
rect 23393 5956 23397 6012
rect 23333 5952 23397 5956
rect 6487 5468 6551 5472
rect 6487 5412 6491 5468
rect 6491 5412 6547 5468
rect 6547 5412 6551 5468
rect 6487 5408 6551 5412
rect 6567 5468 6631 5472
rect 6567 5412 6571 5468
rect 6571 5412 6627 5468
rect 6627 5412 6631 5468
rect 6567 5408 6631 5412
rect 6647 5468 6711 5472
rect 6647 5412 6651 5468
rect 6651 5412 6707 5468
rect 6707 5412 6711 5468
rect 6647 5408 6711 5412
rect 6727 5468 6791 5472
rect 6727 5412 6731 5468
rect 6731 5412 6787 5468
rect 6787 5412 6791 5468
rect 6727 5408 6791 5412
rect 17558 5468 17622 5472
rect 17558 5412 17562 5468
rect 17562 5412 17618 5468
rect 17618 5412 17622 5468
rect 17558 5408 17622 5412
rect 17638 5468 17702 5472
rect 17638 5412 17642 5468
rect 17642 5412 17698 5468
rect 17698 5412 17702 5468
rect 17638 5408 17702 5412
rect 17718 5468 17782 5472
rect 17718 5412 17722 5468
rect 17722 5412 17778 5468
rect 17778 5412 17782 5468
rect 17718 5408 17782 5412
rect 17798 5468 17862 5472
rect 17798 5412 17802 5468
rect 17802 5412 17858 5468
rect 17858 5412 17862 5468
rect 17798 5408 17862 5412
rect 28628 5468 28692 5472
rect 28628 5412 28632 5468
rect 28632 5412 28688 5468
rect 28688 5412 28692 5468
rect 28628 5408 28692 5412
rect 28708 5468 28772 5472
rect 28708 5412 28712 5468
rect 28712 5412 28768 5468
rect 28768 5412 28772 5468
rect 28708 5408 28772 5412
rect 28788 5468 28852 5472
rect 28788 5412 28792 5468
rect 28792 5412 28848 5468
rect 28848 5412 28852 5468
rect 28788 5408 28852 5412
rect 28868 5468 28932 5472
rect 28868 5412 28872 5468
rect 28872 5412 28928 5468
rect 28928 5412 28932 5468
rect 28868 5408 28932 5412
rect 12022 4924 12086 4928
rect 12022 4868 12026 4924
rect 12026 4868 12082 4924
rect 12082 4868 12086 4924
rect 12022 4864 12086 4868
rect 12102 4924 12166 4928
rect 12102 4868 12106 4924
rect 12106 4868 12162 4924
rect 12162 4868 12166 4924
rect 12102 4864 12166 4868
rect 12182 4924 12246 4928
rect 12182 4868 12186 4924
rect 12186 4868 12242 4924
rect 12242 4868 12246 4924
rect 12182 4864 12246 4868
rect 12262 4924 12326 4928
rect 12262 4868 12266 4924
rect 12266 4868 12322 4924
rect 12322 4868 12326 4924
rect 12262 4864 12326 4868
rect 23093 4924 23157 4928
rect 23093 4868 23097 4924
rect 23097 4868 23153 4924
rect 23153 4868 23157 4924
rect 23093 4864 23157 4868
rect 23173 4924 23237 4928
rect 23173 4868 23177 4924
rect 23177 4868 23233 4924
rect 23233 4868 23237 4924
rect 23173 4864 23237 4868
rect 23253 4924 23317 4928
rect 23253 4868 23257 4924
rect 23257 4868 23313 4924
rect 23313 4868 23317 4924
rect 23253 4864 23317 4868
rect 23333 4924 23397 4928
rect 23333 4868 23337 4924
rect 23337 4868 23393 4924
rect 23393 4868 23397 4924
rect 23333 4864 23397 4868
rect 6487 4380 6551 4384
rect 6487 4324 6491 4380
rect 6491 4324 6547 4380
rect 6547 4324 6551 4380
rect 6487 4320 6551 4324
rect 6567 4380 6631 4384
rect 6567 4324 6571 4380
rect 6571 4324 6627 4380
rect 6627 4324 6631 4380
rect 6567 4320 6631 4324
rect 6647 4380 6711 4384
rect 6647 4324 6651 4380
rect 6651 4324 6707 4380
rect 6707 4324 6711 4380
rect 6647 4320 6711 4324
rect 6727 4380 6791 4384
rect 6727 4324 6731 4380
rect 6731 4324 6787 4380
rect 6787 4324 6791 4380
rect 6727 4320 6791 4324
rect 17558 4380 17622 4384
rect 17558 4324 17562 4380
rect 17562 4324 17618 4380
rect 17618 4324 17622 4380
rect 17558 4320 17622 4324
rect 17638 4380 17702 4384
rect 17638 4324 17642 4380
rect 17642 4324 17698 4380
rect 17698 4324 17702 4380
rect 17638 4320 17702 4324
rect 17718 4380 17782 4384
rect 17718 4324 17722 4380
rect 17722 4324 17778 4380
rect 17778 4324 17782 4380
rect 17718 4320 17782 4324
rect 17798 4380 17862 4384
rect 17798 4324 17802 4380
rect 17802 4324 17858 4380
rect 17858 4324 17862 4380
rect 17798 4320 17862 4324
rect 28628 4380 28692 4384
rect 28628 4324 28632 4380
rect 28632 4324 28688 4380
rect 28688 4324 28692 4380
rect 28628 4320 28692 4324
rect 28708 4380 28772 4384
rect 28708 4324 28712 4380
rect 28712 4324 28768 4380
rect 28768 4324 28772 4380
rect 28708 4320 28772 4324
rect 28788 4380 28852 4384
rect 28788 4324 28792 4380
rect 28792 4324 28848 4380
rect 28848 4324 28852 4380
rect 28788 4320 28852 4324
rect 28868 4380 28932 4384
rect 28868 4324 28872 4380
rect 28872 4324 28928 4380
rect 28928 4324 28932 4380
rect 28868 4320 28932 4324
rect 12022 3836 12086 3840
rect 12022 3780 12026 3836
rect 12026 3780 12082 3836
rect 12082 3780 12086 3836
rect 12022 3776 12086 3780
rect 12102 3836 12166 3840
rect 12102 3780 12106 3836
rect 12106 3780 12162 3836
rect 12162 3780 12166 3836
rect 12102 3776 12166 3780
rect 12182 3836 12246 3840
rect 12182 3780 12186 3836
rect 12186 3780 12242 3836
rect 12242 3780 12246 3836
rect 12182 3776 12246 3780
rect 12262 3836 12326 3840
rect 12262 3780 12266 3836
rect 12266 3780 12322 3836
rect 12322 3780 12326 3836
rect 12262 3776 12326 3780
rect 23093 3836 23157 3840
rect 23093 3780 23097 3836
rect 23097 3780 23153 3836
rect 23153 3780 23157 3836
rect 23093 3776 23157 3780
rect 23173 3836 23237 3840
rect 23173 3780 23177 3836
rect 23177 3780 23233 3836
rect 23233 3780 23237 3836
rect 23173 3776 23237 3780
rect 23253 3836 23317 3840
rect 23253 3780 23257 3836
rect 23257 3780 23313 3836
rect 23313 3780 23317 3836
rect 23253 3776 23317 3780
rect 23333 3836 23397 3840
rect 23333 3780 23337 3836
rect 23337 3780 23393 3836
rect 23393 3780 23397 3836
rect 23333 3776 23397 3780
rect 6487 3292 6551 3296
rect 6487 3236 6491 3292
rect 6491 3236 6547 3292
rect 6547 3236 6551 3292
rect 6487 3232 6551 3236
rect 6567 3292 6631 3296
rect 6567 3236 6571 3292
rect 6571 3236 6627 3292
rect 6627 3236 6631 3292
rect 6567 3232 6631 3236
rect 6647 3292 6711 3296
rect 6647 3236 6651 3292
rect 6651 3236 6707 3292
rect 6707 3236 6711 3292
rect 6647 3232 6711 3236
rect 6727 3292 6791 3296
rect 6727 3236 6731 3292
rect 6731 3236 6787 3292
rect 6787 3236 6791 3292
rect 6727 3232 6791 3236
rect 17558 3292 17622 3296
rect 17558 3236 17562 3292
rect 17562 3236 17618 3292
rect 17618 3236 17622 3292
rect 17558 3232 17622 3236
rect 17638 3292 17702 3296
rect 17638 3236 17642 3292
rect 17642 3236 17698 3292
rect 17698 3236 17702 3292
rect 17638 3232 17702 3236
rect 17718 3292 17782 3296
rect 17718 3236 17722 3292
rect 17722 3236 17778 3292
rect 17778 3236 17782 3292
rect 17718 3232 17782 3236
rect 17798 3292 17862 3296
rect 17798 3236 17802 3292
rect 17802 3236 17858 3292
rect 17858 3236 17862 3292
rect 17798 3232 17862 3236
rect 28628 3292 28692 3296
rect 28628 3236 28632 3292
rect 28632 3236 28688 3292
rect 28688 3236 28692 3292
rect 28628 3232 28692 3236
rect 28708 3292 28772 3296
rect 28708 3236 28712 3292
rect 28712 3236 28768 3292
rect 28768 3236 28772 3292
rect 28708 3232 28772 3236
rect 28788 3292 28852 3296
rect 28788 3236 28792 3292
rect 28792 3236 28848 3292
rect 28848 3236 28852 3292
rect 28788 3232 28852 3236
rect 28868 3292 28932 3296
rect 28868 3236 28872 3292
rect 28872 3236 28928 3292
rect 28928 3236 28932 3292
rect 28868 3232 28932 3236
rect 12022 2748 12086 2752
rect 12022 2692 12026 2748
rect 12026 2692 12082 2748
rect 12082 2692 12086 2748
rect 12022 2688 12086 2692
rect 12102 2748 12166 2752
rect 12102 2692 12106 2748
rect 12106 2692 12162 2748
rect 12162 2692 12166 2748
rect 12102 2688 12166 2692
rect 12182 2748 12246 2752
rect 12182 2692 12186 2748
rect 12186 2692 12242 2748
rect 12242 2692 12246 2748
rect 12182 2688 12246 2692
rect 12262 2748 12326 2752
rect 12262 2692 12266 2748
rect 12266 2692 12322 2748
rect 12322 2692 12326 2748
rect 12262 2688 12326 2692
rect 23093 2748 23157 2752
rect 23093 2692 23097 2748
rect 23097 2692 23153 2748
rect 23153 2692 23157 2748
rect 23093 2688 23157 2692
rect 23173 2748 23237 2752
rect 23173 2692 23177 2748
rect 23177 2692 23233 2748
rect 23233 2692 23237 2748
rect 23173 2688 23237 2692
rect 23253 2748 23317 2752
rect 23253 2692 23257 2748
rect 23257 2692 23313 2748
rect 23313 2692 23317 2748
rect 23253 2688 23317 2692
rect 23333 2748 23397 2752
rect 23333 2692 23337 2748
rect 23337 2692 23393 2748
rect 23393 2692 23397 2748
rect 23333 2688 23397 2692
rect 6487 2204 6551 2208
rect 6487 2148 6491 2204
rect 6491 2148 6547 2204
rect 6547 2148 6551 2204
rect 6487 2144 6551 2148
rect 6567 2204 6631 2208
rect 6567 2148 6571 2204
rect 6571 2148 6627 2204
rect 6627 2148 6631 2204
rect 6567 2144 6631 2148
rect 6647 2204 6711 2208
rect 6647 2148 6651 2204
rect 6651 2148 6707 2204
rect 6707 2148 6711 2204
rect 6647 2144 6711 2148
rect 6727 2204 6791 2208
rect 6727 2148 6731 2204
rect 6731 2148 6787 2204
rect 6787 2148 6791 2204
rect 6727 2144 6791 2148
rect 17558 2204 17622 2208
rect 17558 2148 17562 2204
rect 17562 2148 17618 2204
rect 17618 2148 17622 2204
rect 17558 2144 17622 2148
rect 17638 2204 17702 2208
rect 17638 2148 17642 2204
rect 17642 2148 17698 2204
rect 17698 2148 17702 2204
rect 17638 2144 17702 2148
rect 17718 2204 17782 2208
rect 17718 2148 17722 2204
rect 17722 2148 17778 2204
rect 17778 2148 17782 2204
rect 17718 2144 17782 2148
rect 17798 2204 17862 2208
rect 17798 2148 17802 2204
rect 17802 2148 17858 2204
rect 17858 2148 17862 2204
rect 17798 2144 17862 2148
rect 28628 2204 28692 2208
rect 28628 2148 28632 2204
rect 28632 2148 28688 2204
rect 28688 2148 28692 2204
rect 28628 2144 28692 2148
rect 28708 2204 28772 2208
rect 28708 2148 28712 2204
rect 28712 2148 28768 2204
rect 28768 2148 28772 2204
rect 28708 2144 28772 2148
rect 28788 2204 28852 2208
rect 28788 2148 28792 2204
rect 28792 2148 28848 2204
rect 28848 2148 28852 2204
rect 28788 2144 28852 2148
rect 28868 2204 28932 2208
rect 28868 2148 28872 2204
rect 28872 2148 28928 2204
rect 28928 2148 28932 2204
rect 28868 2144 28932 2148
<< metal4 >>
rect 6479 34848 6799 35408
rect 6479 34784 6487 34848
rect 6551 34784 6567 34848
rect 6631 34784 6647 34848
rect 6711 34784 6727 34848
rect 6791 34784 6799 34848
rect 6479 33760 6799 34784
rect 6479 33696 6487 33760
rect 6551 33696 6567 33760
rect 6631 33696 6647 33760
rect 6711 33696 6727 33760
rect 6791 33696 6799 33760
rect 6479 32672 6799 33696
rect 6479 32608 6487 32672
rect 6551 32608 6567 32672
rect 6631 32608 6647 32672
rect 6711 32608 6727 32672
rect 6791 32608 6799 32672
rect 6479 31584 6799 32608
rect 6479 31520 6487 31584
rect 6551 31520 6567 31584
rect 6631 31520 6647 31584
rect 6711 31520 6727 31584
rect 6791 31520 6799 31584
rect 6479 30496 6799 31520
rect 6479 30432 6487 30496
rect 6551 30432 6567 30496
rect 6631 30432 6647 30496
rect 6711 30432 6727 30496
rect 6791 30432 6799 30496
rect 6479 29899 6799 30432
rect 6479 29663 6521 29899
rect 6757 29663 6799 29899
rect 6479 29408 6799 29663
rect 6479 29344 6487 29408
rect 6551 29344 6567 29408
rect 6631 29344 6647 29408
rect 6711 29344 6727 29408
rect 6791 29344 6799 29408
rect 6479 28320 6799 29344
rect 6479 28256 6487 28320
rect 6551 28256 6567 28320
rect 6631 28256 6647 28320
rect 6711 28256 6727 28320
rect 6791 28256 6799 28320
rect 6479 27232 6799 28256
rect 6479 27168 6487 27232
rect 6551 27168 6567 27232
rect 6631 27168 6647 27232
rect 6711 27168 6727 27232
rect 6791 27168 6799 27232
rect 6479 26144 6799 27168
rect 6479 26080 6487 26144
rect 6551 26080 6567 26144
rect 6631 26080 6647 26144
rect 6711 26080 6727 26144
rect 6791 26080 6799 26144
rect 6479 25056 6799 26080
rect 6479 24992 6487 25056
rect 6551 24992 6567 25056
rect 6631 24992 6647 25056
rect 6711 24992 6727 25056
rect 6791 24992 6799 25056
rect 6479 23968 6799 24992
rect 6479 23904 6487 23968
rect 6551 23904 6567 23968
rect 6631 23904 6647 23968
rect 6711 23904 6727 23968
rect 6791 23904 6799 23968
rect 6479 22880 6799 23904
rect 6479 22816 6487 22880
rect 6551 22816 6567 22880
rect 6631 22816 6647 22880
rect 6711 22816 6727 22880
rect 6791 22816 6799 22880
rect 6479 21792 6799 22816
rect 6479 21728 6487 21792
rect 6551 21728 6567 21792
rect 6631 21728 6647 21792
rect 6711 21728 6727 21792
rect 6791 21728 6799 21792
rect 6479 20704 6799 21728
rect 6479 20640 6487 20704
rect 6551 20640 6567 20704
rect 6631 20640 6647 20704
rect 6711 20640 6727 20704
rect 6791 20640 6799 20704
rect 6479 19616 6799 20640
rect 6479 19552 6487 19616
rect 6551 19552 6567 19616
rect 6631 19552 6647 19616
rect 6711 19552 6727 19616
rect 6791 19552 6799 19616
rect 6479 18838 6799 19552
rect 6479 18602 6521 18838
rect 6757 18602 6799 18838
rect 6479 18528 6799 18602
rect 6479 18464 6487 18528
rect 6551 18464 6567 18528
rect 6631 18464 6647 18528
rect 6711 18464 6727 18528
rect 6791 18464 6799 18528
rect 6479 17440 6799 18464
rect 6479 17376 6487 17440
rect 6551 17376 6567 17440
rect 6631 17376 6647 17440
rect 6711 17376 6727 17440
rect 6791 17376 6799 17440
rect 6479 16352 6799 17376
rect 6479 16288 6487 16352
rect 6551 16288 6567 16352
rect 6631 16288 6647 16352
rect 6711 16288 6727 16352
rect 6791 16288 6799 16352
rect 6479 15264 6799 16288
rect 6479 15200 6487 15264
rect 6551 15200 6567 15264
rect 6631 15200 6647 15264
rect 6711 15200 6727 15264
rect 6791 15200 6799 15264
rect 6479 14176 6799 15200
rect 6479 14112 6487 14176
rect 6551 14112 6567 14176
rect 6631 14112 6647 14176
rect 6711 14112 6727 14176
rect 6791 14112 6799 14176
rect 6479 13088 6799 14112
rect 6479 13024 6487 13088
rect 6551 13024 6567 13088
rect 6631 13024 6647 13088
rect 6711 13024 6727 13088
rect 6791 13024 6799 13088
rect 6479 12000 6799 13024
rect 6479 11936 6487 12000
rect 6551 11936 6567 12000
rect 6631 11936 6647 12000
rect 6711 11936 6727 12000
rect 6791 11936 6799 12000
rect 6479 10912 6799 11936
rect 6479 10848 6487 10912
rect 6551 10848 6567 10912
rect 6631 10848 6647 10912
rect 6711 10848 6727 10912
rect 6791 10848 6799 10912
rect 6479 9824 6799 10848
rect 6479 9760 6487 9824
rect 6551 9760 6567 9824
rect 6631 9760 6647 9824
rect 6711 9760 6727 9824
rect 6791 9760 6799 9824
rect 6479 8736 6799 9760
rect 6479 8672 6487 8736
rect 6551 8672 6567 8736
rect 6631 8672 6647 8736
rect 6711 8672 6727 8736
rect 6791 8672 6799 8736
rect 6479 7776 6799 8672
rect 6479 7648 6521 7776
rect 6757 7648 6799 7776
rect 6479 7584 6487 7648
rect 6791 7584 6799 7648
rect 6479 7540 6521 7584
rect 6757 7540 6799 7584
rect 6479 6560 6799 7540
rect 6479 6496 6487 6560
rect 6551 6496 6567 6560
rect 6631 6496 6647 6560
rect 6711 6496 6727 6560
rect 6791 6496 6799 6560
rect 6479 5472 6799 6496
rect 6479 5408 6487 5472
rect 6551 5408 6567 5472
rect 6631 5408 6647 5472
rect 6711 5408 6727 5472
rect 6791 5408 6799 5472
rect 6479 4384 6799 5408
rect 6479 4320 6487 4384
rect 6551 4320 6567 4384
rect 6631 4320 6647 4384
rect 6711 4320 6727 4384
rect 6791 4320 6799 4384
rect 6479 3296 6799 4320
rect 6479 3232 6487 3296
rect 6551 3232 6567 3296
rect 6631 3232 6647 3296
rect 6711 3232 6727 3296
rect 6791 3232 6799 3296
rect 6479 2208 6799 3232
rect 6479 2144 6487 2208
rect 6551 2144 6567 2208
rect 6631 2144 6647 2208
rect 6711 2144 6727 2208
rect 6791 2144 6799 2208
rect 6479 2128 6799 2144
rect 12014 35392 12335 35408
rect 12014 35328 12022 35392
rect 12086 35328 12102 35392
rect 12166 35328 12182 35392
rect 12246 35328 12262 35392
rect 12326 35328 12335 35392
rect 12014 34304 12335 35328
rect 12014 34240 12022 34304
rect 12086 34240 12102 34304
rect 12166 34240 12182 34304
rect 12246 34240 12262 34304
rect 12326 34240 12335 34304
rect 12014 33216 12335 34240
rect 12014 33152 12022 33216
rect 12086 33152 12102 33216
rect 12166 33152 12182 33216
rect 12246 33152 12262 33216
rect 12326 33152 12335 33216
rect 12014 32128 12335 33152
rect 12014 32064 12022 32128
rect 12086 32064 12102 32128
rect 12166 32064 12182 32128
rect 12246 32064 12262 32128
rect 12326 32064 12335 32128
rect 12014 31040 12335 32064
rect 12014 30976 12022 31040
rect 12086 30976 12102 31040
rect 12166 30976 12182 31040
rect 12246 30976 12262 31040
rect 12326 30976 12335 31040
rect 12014 29952 12335 30976
rect 12014 29888 12022 29952
rect 12086 29888 12102 29952
rect 12166 29888 12182 29952
rect 12246 29888 12262 29952
rect 12326 29888 12335 29952
rect 12014 28864 12335 29888
rect 12014 28800 12022 28864
rect 12086 28800 12102 28864
rect 12166 28800 12182 28864
rect 12246 28800 12262 28864
rect 12326 28800 12335 28864
rect 12014 27776 12335 28800
rect 12014 27712 12022 27776
rect 12086 27712 12102 27776
rect 12166 27712 12182 27776
rect 12246 27712 12262 27776
rect 12326 27712 12335 27776
rect 12014 26688 12335 27712
rect 12014 26624 12022 26688
rect 12086 26624 12102 26688
rect 12166 26624 12182 26688
rect 12246 26624 12262 26688
rect 12326 26624 12335 26688
rect 12014 25600 12335 26624
rect 12014 25536 12022 25600
rect 12086 25536 12102 25600
rect 12166 25536 12182 25600
rect 12246 25536 12262 25600
rect 12326 25536 12335 25600
rect 12014 24512 12335 25536
rect 12014 24448 12022 24512
rect 12086 24448 12102 24512
rect 12166 24448 12182 24512
rect 12246 24448 12262 24512
rect 12326 24448 12335 24512
rect 12014 24368 12335 24448
rect 12014 24132 12056 24368
rect 12292 24132 12335 24368
rect 12014 23424 12335 24132
rect 12014 23360 12022 23424
rect 12086 23360 12102 23424
rect 12166 23360 12182 23424
rect 12246 23360 12262 23424
rect 12326 23360 12335 23424
rect 12014 22336 12335 23360
rect 12014 22272 12022 22336
rect 12086 22272 12102 22336
rect 12166 22272 12182 22336
rect 12246 22272 12262 22336
rect 12326 22272 12335 22336
rect 12014 21248 12335 22272
rect 12014 21184 12022 21248
rect 12086 21184 12102 21248
rect 12166 21184 12182 21248
rect 12246 21184 12262 21248
rect 12326 21184 12335 21248
rect 12014 20160 12335 21184
rect 12014 20096 12022 20160
rect 12086 20096 12102 20160
rect 12166 20096 12182 20160
rect 12246 20096 12262 20160
rect 12326 20096 12335 20160
rect 12014 19072 12335 20096
rect 12014 19008 12022 19072
rect 12086 19008 12102 19072
rect 12166 19008 12182 19072
rect 12246 19008 12262 19072
rect 12326 19008 12335 19072
rect 12014 17984 12335 19008
rect 12014 17920 12022 17984
rect 12086 17920 12102 17984
rect 12166 17920 12182 17984
rect 12246 17920 12262 17984
rect 12326 17920 12335 17984
rect 12014 16896 12335 17920
rect 12014 16832 12022 16896
rect 12086 16832 12102 16896
rect 12166 16832 12182 16896
rect 12246 16832 12262 16896
rect 12326 16832 12335 16896
rect 12014 15808 12335 16832
rect 12014 15744 12022 15808
rect 12086 15744 12102 15808
rect 12166 15744 12182 15808
rect 12246 15744 12262 15808
rect 12326 15744 12335 15808
rect 12014 14720 12335 15744
rect 12014 14656 12022 14720
rect 12086 14656 12102 14720
rect 12166 14656 12182 14720
rect 12246 14656 12262 14720
rect 12326 14656 12335 14720
rect 12014 13632 12335 14656
rect 12014 13568 12022 13632
rect 12086 13568 12102 13632
rect 12166 13568 12182 13632
rect 12246 13568 12262 13632
rect 12326 13568 12335 13632
rect 12014 13307 12335 13568
rect 12014 13071 12056 13307
rect 12292 13071 12335 13307
rect 12014 12544 12335 13071
rect 12014 12480 12022 12544
rect 12086 12480 12102 12544
rect 12166 12480 12182 12544
rect 12246 12480 12262 12544
rect 12326 12480 12335 12544
rect 12014 11456 12335 12480
rect 12014 11392 12022 11456
rect 12086 11392 12102 11456
rect 12166 11392 12182 11456
rect 12246 11392 12262 11456
rect 12326 11392 12335 11456
rect 12014 10368 12335 11392
rect 12014 10304 12022 10368
rect 12086 10304 12102 10368
rect 12166 10304 12182 10368
rect 12246 10304 12262 10368
rect 12326 10304 12335 10368
rect 12014 9280 12335 10304
rect 12014 9216 12022 9280
rect 12086 9216 12102 9280
rect 12166 9216 12182 9280
rect 12246 9216 12262 9280
rect 12326 9216 12335 9280
rect 12014 8192 12335 9216
rect 12014 8128 12022 8192
rect 12086 8128 12102 8192
rect 12166 8128 12182 8192
rect 12246 8128 12262 8192
rect 12326 8128 12335 8192
rect 12014 7104 12335 8128
rect 12014 7040 12022 7104
rect 12086 7040 12102 7104
rect 12166 7040 12182 7104
rect 12246 7040 12262 7104
rect 12326 7040 12335 7104
rect 12014 6016 12335 7040
rect 12014 5952 12022 6016
rect 12086 5952 12102 6016
rect 12166 5952 12182 6016
rect 12246 5952 12262 6016
rect 12326 5952 12335 6016
rect 12014 4928 12335 5952
rect 12014 4864 12022 4928
rect 12086 4864 12102 4928
rect 12166 4864 12182 4928
rect 12246 4864 12262 4928
rect 12326 4864 12335 4928
rect 12014 3840 12335 4864
rect 12014 3776 12022 3840
rect 12086 3776 12102 3840
rect 12166 3776 12182 3840
rect 12246 3776 12262 3840
rect 12326 3776 12335 3840
rect 12014 2752 12335 3776
rect 12014 2688 12022 2752
rect 12086 2688 12102 2752
rect 12166 2688 12182 2752
rect 12246 2688 12262 2752
rect 12326 2688 12335 2752
rect 12014 2128 12335 2688
rect 17550 34848 17870 35408
rect 17550 34784 17558 34848
rect 17622 34784 17638 34848
rect 17702 34784 17718 34848
rect 17782 34784 17798 34848
rect 17862 34784 17870 34848
rect 17550 33760 17870 34784
rect 17550 33696 17558 33760
rect 17622 33696 17638 33760
rect 17702 33696 17718 33760
rect 17782 33696 17798 33760
rect 17862 33696 17870 33760
rect 17550 32672 17870 33696
rect 17550 32608 17558 32672
rect 17622 32608 17638 32672
rect 17702 32608 17718 32672
rect 17782 32608 17798 32672
rect 17862 32608 17870 32672
rect 17550 31584 17870 32608
rect 17550 31520 17558 31584
rect 17622 31520 17638 31584
rect 17702 31520 17718 31584
rect 17782 31520 17798 31584
rect 17862 31520 17870 31584
rect 17550 30496 17870 31520
rect 17550 30432 17558 30496
rect 17622 30432 17638 30496
rect 17702 30432 17718 30496
rect 17782 30432 17798 30496
rect 17862 30432 17870 30496
rect 17550 29899 17870 30432
rect 17550 29663 17592 29899
rect 17828 29663 17870 29899
rect 17550 29408 17870 29663
rect 17550 29344 17558 29408
rect 17622 29344 17638 29408
rect 17702 29344 17718 29408
rect 17782 29344 17798 29408
rect 17862 29344 17870 29408
rect 17550 28320 17870 29344
rect 17550 28256 17558 28320
rect 17622 28256 17638 28320
rect 17702 28256 17718 28320
rect 17782 28256 17798 28320
rect 17862 28256 17870 28320
rect 17550 27232 17870 28256
rect 17550 27168 17558 27232
rect 17622 27168 17638 27232
rect 17702 27168 17718 27232
rect 17782 27168 17798 27232
rect 17862 27168 17870 27232
rect 17550 26144 17870 27168
rect 17550 26080 17558 26144
rect 17622 26080 17638 26144
rect 17702 26080 17718 26144
rect 17782 26080 17798 26144
rect 17862 26080 17870 26144
rect 17550 25056 17870 26080
rect 17550 24992 17558 25056
rect 17622 24992 17638 25056
rect 17702 24992 17718 25056
rect 17782 24992 17798 25056
rect 17862 24992 17870 25056
rect 17550 23968 17870 24992
rect 17550 23904 17558 23968
rect 17622 23904 17638 23968
rect 17702 23904 17718 23968
rect 17782 23904 17798 23968
rect 17862 23904 17870 23968
rect 17550 22880 17870 23904
rect 17550 22816 17558 22880
rect 17622 22816 17638 22880
rect 17702 22816 17718 22880
rect 17782 22816 17798 22880
rect 17862 22816 17870 22880
rect 17550 21792 17870 22816
rect 17550 21728 17558 21792
rect 17622 21728 17638 21792
rect 17702 21728 17718 21792
rect 17782 21728 17798 21792
rect 17862 21728 17870 21792
rect 17550 20704 17870 21728
rect 17550 20640 17558 20704
rect 17622 20640 17638 20704
rect 17702 20640 17718 20704
rect 17782 20640 17798 20704
rect 17862 20640 17870 20704
rect 17550 19616 17870 20640
rect 17550 19552 17558 19616
rect 17622 19552 17638 19616
rect 17702 19552 17718 19616
rect 17782 19552 17798 19616
rect 17862 19552 17870 19616
rect 17550 18838 17870 19552
rect 17550 18602 17592 18838
rect 17828 18602 17870 18838
rect 17550 18528 17870 18602
rect 17550 18464 17558 18528
rect 17622 18464 17638 18528
rect 17702 18464 17718 18528
rect 17782 18464 17798 18528
rect 17862 18464 17870 18528
rect 17550 17440 17870 18464
rect 17550 17376 17558 17440
rect 17622 17376 17638 17440
rect 17702 17376 17718 17440
rect 17782 17376 17798 17440
rect 17862 17376 17870 17440
rect 17550 16352 17870 17376
rect 17550 16288 17558 16352
rect 17622 16288 17638 16352
rect 17702 16288 17718 16352
rect 17782 16288 17798 16352
rect 17862 16288 17870 16352
rect 17550 15264 17870 16288
rect 17550 15200 17558 15264
rect 17622 15200 17638 15264
rect 17702 15200 17718 15264
rect 17782 15200 17798 15264
rect 17862 15200 17870 15264
rect 17550 14176 17870 15200
rect 17550 14112 17558 14176
rect 17622 14112 17638 14176
rect 17702 14112 17718 14176
rect 17782 14112 17798 14176
rect 17862 14112 17870 14176
rect 17550 13088 17870 14112
rect 17550 13024 17558 13088
rect 17622 13024 17638 13088
rect 17702 13024 17718 13088
rect 17782 13024 17798 13088
rect 17862 13024 17870 13088
rect 17550 12000 17870 13024
rect 17550 11936 17558 12000
rect 17622 11936 17638 12000
rect 17702 11936 17718 12000
rect 17782 11936 17798 12000
rect 17862 11936 17870 12000
rect 17550 10912 17870 11936
rect 17550 10848 17558 10912
rect 17622 10848 17638 10912
rect 17702 10848 17718 10912
rect 17782 10848 17798 10912
rect 17862 10848 17870 10912
rect 17550 9824 17870 10848
rect 17550 9760 17558 9824
rect 17622 9760 17638 9824
rect 17702 9760 17718 9824
rect 17782 9760 17798 9824
rect 17862 9760 17870 9824
rect 17550 8736 17870 9760
rect 17550 8672 17558 8736
rect 17622 8672 17638 8736
rect 17702 8672 17718 8736
rect 17782 8672 17798 8736
rect 17862 8672 17870 8736
rect 17550 7776 17870 8672
rect 17550 7648 17592 7776
rect 17828 7648 17870 7776
rect 17550 7584 17558 7648
rect 17862 7584 17870 7648
rect 17550 7540 17592 7584
rect 17828 7540 17870 7584
rect 17550 6560 17870 7540
rect 17550 6496 17558 6560
rect 17622 6496 17638 6560
rect 17702 6496 17718 6560
rect 17782 6496 17798 6560
rect 17862 6496 17870 6560
rect 17550 5472 17870 6496
rect 17550 5408 17558 5472
rect 17622 5408 17638 5472
rect 17702 5408 17718 5472
rect 17782 5408 17798 5472
rect 17862 5408 17870 5472
rect 17550 4384 17870 5408
rect 17550 4320 17558 4384
rect 17622 4320 17638 4384
rect 17702 4320 17718 4384
rect 17782 4320 17798 4384
rect 17862 4320 17870 4384
rect 17550 3296 17870 4320
rect 17550 3232 17558 3296
rect 17622 3232 17638 3296
rect 17702 3232 17718 3296
rect 17782 3232 17798 3296
rect 17862 3232 17870 3296
rect 17550 2208 17870 3232
rect 17550 2144 17558 2208
rect 17622 2144 17638 2208
rect 17702 2144 17718 2208
rect 17782 2144 17798 2208
rect 17862 2144 17870 2208
rect 17550 2128 17870 2144
rect 23085 35392 23405 35408
rect 23085 35328 23093 35392
rect 23157 35328 23173 35392
rect 23237 35328 23253 35392
rect 23317 35328 23333 35392
rect 23397 35328 23405 35392
rect 23085 34304 23405 35328
rect 23085 34240 23093 34304
rect 23157 34240 23173 34304
rect 23237 34240 23253 34304
rect 23317 34240 23333 34304
rect 23397 34240 23405 34304
rect 23085 33216 23405 34240
rect 23085 33152 23093 33216
rect 23157 33152 23173 33216
rect 23237 33152 23253 33216
rect 23317 33152 23333 33216
rect 23397 33152 23405 33216
rect 23085 32128 23405 33152
rect 23085 32064 23093 32128
rect 23157 32064 23173 32128
rect 23237 32064 23253 32128
rect 23317 32064 23333 32128
rect 23397 32064 23405 32128
rect 23085 31040 23405 32064
rect 23085 30976 23093 31040
rect 23157 30976 23173 31040
rect 23237 30976 23253 31040
rect 23317 30976 23333 31040
rect 23397 30976 23405 31040
rect 23085 29952 23405 30976
rect 23085 29888 23093 29952
rect 23157 29888 23173 29952
rect 23237 29888 23253 29952
rect 23317 29888 23333 29952
rect 23397 29888 23405 29952
rect 23085 28864 23405 29888
rect 23085 28800 23093 28864
rect 23157 28800 23173 28864
rect 23237 28800 23253 28864
rect 23317 28800 23333 28864
rect 23397 28800 23405 28864
rect 23085 27776 23405 28800
rect 23085 27712 23093 27776
rect 23157 27712 23173 27776
rect 23237 27712 23253 27776
rect 23317 27712 23333 27776
rect 23397 27712 23405 27776
rect 23085 26688 23405 27712
rect 23085 26624 23093 26688
rect 23157 26624 23173 26688
rect 23237 26624 23253 26688
rect 23317 26624 23333 26688
rect 23397 26624 23405 26688
rect 23085 25600 23405 26624
rect 23085 25536 23093 25600
rect 23157 25536 23173 25600
rect 23237 25536 23253 25600
rect 23317 25536 23333 25600
rect 23397 25536 23405 25600
rect 23085 24512 23405 25536
rect 23085 24448 23093 24512
rect 23157 24448 23173 24512
rect 23237 24448 23253 24512
rect 23317 24448 23333 24512
rect 23397 24448 23405 24512
rect 23085 24368 23405 24448
rect 23085 24132 23127 24368
rect 23363 24132 23405 24368
rect 23085 23424 23405 24132
rect 23085 23360 23093 23424
rect 23157 23360 23173 23424
rect 23237 23360 23253 23424
rect 23317 23360 23333 23424
rect 23397 23360 23405 23424
rect 23085 22336 23405 23360
rect 23085 22272 23093 22336
rect 23157 22272 23173 22336
rect 23237 22272 23253 22336
rect 23317 22272 23333 22336
rect 23397 22272 23405 22336
rect 23085 21248 23405 22272
rect 23085 21184 23093 21248
rect 23157 21184 23173 21248
rect 23237 21184 23253 21248
rect 23317 21184 23333 21248
rect 23397 21184 23405 21248
rect 23085 20160 23405 21184
rect 23085 20096 23093 20160
rect 23157 20096 23173 20160
rect 23237 20096 23253 20160
rect 23317 20096 23333 20160
rect 23397 20096 23405 20160
rect 23085 19072 23405 20096
rect 23085 19008 23093 19072
rect 23157 19008 23173 19072
rect 23237 19008 23253 19072
rect 23317 19008 23333 19072
rect 23397 19008 23405 19072
rect 23085 17984 23405 19008
rect 23085 17920 23093 17984
rect 23157 17920 23173 17984
rect 23237 17920 23253 17984
rect 23317 17920 23333 17984
rect 23397 17920 23405 17984
rect 23085 16896 23405 17920
rect 23085 16832 23093 16896
rect 23157 16832 23173 16896
rect 23237 16832 23253 16896
rect 23317 16832 23333 16896
rect 23397 16832 23405 16896
rect 23085 15808 23405 16832
rect 23085 15744 23093 15808
rect 23157 15744 23173 15808
rect 23237 15744 23253 15808
rect 23317 15744 23333 15808
rect 23397 15744 23405 15808
rect 23085 14720 23405 15744
rect 23085 14656 23093 14720
rect 23157 14656 23173 14720
rect 23237 14656 23253 14720
rect 23317 14656 23333 14720
rect 23397 14656 23405 14720
rect 23085 13632 23405 14656
rect 23085 13568 23093 13632
rect 23157 13568 23173 13632
rect 23237 13568 23253 13632
rect 23317 13568 23333 13632
rect 23397 13568 23405 13632
rect 23085 13307 23405 13568
rect 23085 13071 23127 13307
rect 23363 13071 23405 13307
rect 23085 12544 23405 13071
rect 23085 12480 23093 12544
rect 23157 12480 23173 12544
rect 23237 12480 23253 12544
rect 23317 12480 23333 12544
rect 23397 12480 23405 12544
rect 23085 11456 23405 12480
rect 23085 11392 23093 11456
rect 23157 11392 23173 11456
rect 23237 11392 23253 11456
rect 23317 11392 23333 11456
rect 23397 11392 23405 11456
rect 23085 10368 23405 11392
rect 23085 10304 23093 10368
rect 23157 10304 23173 10368
rect 23237 10304 23253 10368
rect 23317 10304 23333 10368
rect 23397 10304 23405 10368
rect 23085 9280 23405 10304
rect 23085 9216 23093 9280
rect 23157 9216 23173 9280
rect 23237 9216 23253 9280
rect 23317 9216 23333 9280
rect 23397 9216 23405 9280
rect 23085 8192 23405 9216
rect 23085 8128 23093 8192
rect 23157 8128 23173 8192
rect 23237 8128 23253 8192
rect 23317 8128 23333 8192
rect 23397 8128 23405 8192
rect 23085 7104 23405 8128
rect 23085 7040 23093 7104
rect 23157 7040 23173 7104
rect 23237 7040 23253 7104
rect 23317 7040 23333 7104
rect 23397 7040 23405 7104
rect 23085 6016 23405 7040
rect 23085 5952 23093 6016
rect 23157 5952 23173 6016
rect 23237 5952 23253 6016
rect 23317 5952 23333 6016
rect 23397 5952 23405 6016
rect 23085 4928 23405 5952
rect 23085 4864 23093 4928
rect 23157 4864 23173 4928
rect 23237 4864 23253 4928
rect 23317 4864 23333 4928
rect 23397 4864 23405 4928
rect 23085 3840 23405 4864
rect 23085 3776 23093 3840
rect 23157 3776 23173 3840
rect 23237 3776 23253 3840
rect 23317 3776 23333 3840
rect 23397 3776 23405 3840
rect 23085 2752 23405 3776
rect 23085 2688 23093 2752
rect 23157 2688 23173 2752
rect 23237 2688 23253 2752
rect 23317 2688 23333 2752
rect 23397 2688 23405 2752
rect 23085 2128 23405 2688
rect 28620 34848 28941 35408
rect 28620 34784 28628 34848
rect 28692 34784 28708 34848
rect 28772 34784 28788 34848
rect 28852 34784 28868 34848
rect 28932 34784 28941 34848
rect 28620 33760 28941 34784
rect 28620 33696 28628 33760
rect 28692 33696 28708 33760
rect 28772 33696 28788 33760
rect 28852 33696 28868 33760
rect 28932 33696 28941 33760
rect 28620 32672 28941 33696
rect 28620 32608 28628 32672
rect 28692 32608 28708 32672
rect 28772 32608 28788 32672
rect 28852 32608 28868 32672
rect 28932 32608 28941 32672
rect 28620 31584 28941 32608
rect 28620 31520 28628 31584
rect 28692 31520 28708 31584
rect 28772 31520 28788 31584
rect 28852 31520 28868 31584
rect 28932 31520 28941 31584
rect 28620 30496 28941 31520
rect 28620 30432 28628 30496
rect 28692 30432 28708 30496
rect 28772 30432 28788 30496
rect 28852 30432 28868 30496
rect 28932 30432 28941 30496
rect 28620 29899 28941 30432
rect 28620 29663 28662 29899
rect 28898 29663 28941 29899
rect 28620 29408 28941 29663
rect 28620 29344 28628 29408
rect 28692 29344 28708 29408
rect 28772 29344 28788 29408
rect 28852 29344 28868 29408
rect 28932 29344 28941 29408
rect 28620 28320 28941 29344
rect 28620 28256 28628 28320
rect 28692 28256 28708 28320
rect 28772 28256 28788 28320
rect 28852 28256 28868 28320
rect 28932 28256 28941 28320
rect 28620 27232 28941 28256
rect 28620 27168 28628 27232
rect 28692 27168 28708 27232
rect 28772 27168 28788 27232
rect 28852 27168 28868 27232
rect 28932 27168 28941 27232
rect 28620 26144 28941 27168
rect 28620 26080 28628 26144
rect 28692 26080 28708 26144
rect 28772 26080 28788 26144
rect 28852 26080 28868 26144
rect 28932 26080 28941 26144
rect 28620 25056 28941 26080
rect 28620 24992 28628 25056
rect 28692 24992 28708 25056
rect 28772 24992 28788 25056
rect 28852 24992 28868 25056
rect 28932 24992 28941 25056
rect 28620 23968 28941 24992
rect 28620 23904 28628 23968
rect 28692 23904 28708 23968
rect 28772 23904 28788 23968
rect 28852 23904 28868 23968
rect 28932 23904 28941 23968
rect 28620 22880 28941 23904
rect 28620 22816 28628 22880
rect 28692 22816 28708 22880
rect 28772 22816 28788 22880
rect 28852 22816 28868 22880
rect 28932 22816 28941 22880
rect 28620 21792 28941 22816
rect 28620 21728 28628 21792
rect 28692 21728 28708 21792
rect 28772 21728 28788 21792
rect 28852 21728 28868 21792
rect 28932 21728 28941 21792
rect 28620 20704 28941 21728
rect 28620 20640 28628 20704
rect 28692 20640 28708 20704
rect 28772 20640 28788 20704
rect 28852 20640 28868 20704
rect 28932 20640 28941 20704
rect 28620 19616 28941 20640
rect 28620 19552 28628 19616
rect 28692 19552 28708 19616
rect 28772 19552 28788 19616
rect 28852 19552 28868 19616
rect 28932 19552 28941 19616
rect 28620 18838 28941 19552
rect 28620 18602 28662 18838
rect 28898 18602 28941 18838
rect 28620 18528 28941 18602
rect 28620 18464 28628 18528
rect 28692 18464 28708 18528
rect 28772 18464 28788 18528
rect 28852 18464 28868 18528
rect 28932 18464 28941 18528
rect 28620 17440 28941 18464
rect 28620 17376 28628 17440
rect 28692 17376 28708 17440
rect 28772 17376 28788 17440
rect 28852 17376 28868 17440
rect 28932 17376 28941 17440
rect 28620 16352 28941 17376
rect 28620 16288 28628 16352
rect 28692 16288 28708 16352
rect 28772 16288 28788 16352
rect 28852 16288 28868 16352
rect 28932 16288 28941 16352
rect 28620 15264 28941 16288
rect 28620 15200 28628 15264
rect 28692 15200 28708 15264
rect 28772 15200 28788 15264
rect 28852 15200 28868 15264
rect 28932 15200 28941 15264
rect 28620 14176 28941 15200
rect 28620 14112 28628 14176
rect 28692 14112 28708 14176
rect 28772 14112 28788 14176
rect 28852 14112 28868 14176
rect 28932 14112 28941 14176
rect 28620 13088 28941 14112
rect 28620 13024 28628 13088
rect 28692 13024 28708 13088
rect 28772 13024 28788 13088
rect 28852 13024 28868 13088
rect 28932 13024 28941 13088
rect 28620 12000 28941 13024
rect 28620 11936 28628 12000
rect 28692 11936 28708 12000
rect 28772 11936 28788 12000
rect 28852 11936 28868 12000
rect 28932 11936 28941 12000
rect 28620 10912 28941 11936
rect 28620 10848 28628 10912
rect 28692 10848 28708 10912
rect 28772 10848 28788 10912
rect 28852 10848 28868 10912
rect 28932 10848 28941 10912
rect 28620 9824 28941 10848
rect 28620 9760 28628 9824
rect 28692 9760 28708 9824
rect 28772 9760 28788 9824
rect 28852 9760 28868 9824
rect 28932 9760 28941 9824
rect 28620 8736 28941 9760
rect 28620 8672 28628 8736
rect 28692 8672 28708 8736
rect 28772 8672 28788 8736
rect 28852 8672 28868 8736
rect 28932 8672 28941 8736
rect 28620 7776 28941 8672
rect 28620 7648 28662 7776
rect 28898 7648 28941 7776
rect 28620 7584 28628 7648
rect 28932 7584 28941 7648
rect 28620 7540 28662 7584
rect 28898 7540 28941 7584
rect 28620 6560 28941 7540
rect 28620 6496 28628 6560
rect 28692 6496 28708 6560
rect 28772 6496 28788 6560
rect 28852 6496 28868 6560
rect 28932 6496 28941 6560
rect 28620 5472 28941 6496
rect 28620 5408 28628 5472
rect 28692 5408 28708 5472
rect 28772 5408 28788 5472
rect 28852 5408 28868 5472
rect 28932 5408 28941 5472
rect 28620 4384 28941 5408
rect 28620 4320 28628 4384
rect 28692 4320 28708 4384
rect 28772 4320 28788 4384
rect 28852 4320 28868 4384
rect 28932 4320 28941 4384
rect 28620 3296 28941 4320
rect 28620 3232 28628 3296
rect 28692 3232 28708 3296
rect 28772 3232 28788 3296
rect 28852 3232 28868 3296
rect 28932 3232 28941 3296
rect 28620 2208 28941 3232
rect 28620 2144 28628 2208
rect 28692 2144 28708 2208
rect 28772 2144 28788 2208
rect 28852 2144 28868 2208
rect 28932 2144 28941 2208
rect 28620 2128 28941 2144
<< via4 >>
rect 6521 29663 6757 29899
rect 6521 18602 6757 18838
rect 6521 7648 6757 7776
rect 6521 7584 6551 7648
rect 6551 7584 6567 7648
rect 6567 7584 6631 7648
rect 6631 7584 6647 7648
rect 6647 7584 6711 7648
rect 6711 7584 6727 7648
rect 6727 7584 6757 7648
rect 6521 7540 6757 7584
rect 12056 24132 12292 24368
rect 12056 13071 12292 13307
rect 17592 29663 17828 29899
rect 17592 18602 17828 18838
rect 17592 7648 17828 7776
rect 17592 7584 17622 7648
rect 17622 7584 17638 7648
rect 17638 7584 17702 7648
rect 17702 7584 17718 7648
rect 17718 7584 17782 7648
rect 17782 7584 17798 7648
rect 17798 7584 17828 7648
rect 17592 7540 17828 7584
rect 23127 24132 23363 24368
rect 23127 13071 23363 13307
rect 28662 29663 28898 29899
rect 28662 18602 28898 18838
rect 28662 7648 28898 7776
rect 28662 7584 28692 7648
rect 28692 7584 28708 7648
rect 28708 7584 28772 7648
rect 28772 7584 28788 7648
rect 28788 7584 28852 7648
rect 28852 7584 28868 7648
rect 28868 7584 28898 7648
rect 28662 7540 28898 7584
<< metal5 >>
rect 1104 29899 34316 29941
rect 1104 29663 6521 29899
rect 6757 29663 17592 29899
rect 17828 29663 28662 29899
rect 28898 29663 34316 29899
rect 1104 29621 34316 29663
rect 1104 24368 34316 24411
rect 1104 24132 12056 24368
rect 12292 24132 23127 24368
rect 23363 24132 34316 24368
rect 1104 24090 34316 24132
rect 1104 18838 34316 18880
rect 1104 18602 6521 18838
rect 6757 18602 17592 18838
rect 17828 18602 28662 18838
rect 28898 18602 34316 18838
rect 1104 18560 34316 18602
rect 1104 13307 34316 13349
rect 1104 13071 12056 13307
rect 12292 13071 23127 13307
rect 23363 13071 34316 13307
rect 1104 13029 34316 13071
rect 1104 7776 34316 7819
rect 1104 7540 6521 7776
rect 6757 7540 17592 7776
rect 17828 7540 28662 7776
rect 28898 7540 34316 7776
rect 1104 7498 34316 7540
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1738175533
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1738175533
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output32
timestamp 1738175533
transform -1 0 2116 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3
timestamp 1738175533
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11
timestamp 1738175533
transform 1 0 2116 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1738175533
transform 1 0 2760 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17
timestamp 1738175533
transform 1 0 2668 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22
timestamp 1738175533
transform 1 0 3128 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1738175533
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1738175533
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1738175533
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28
timestamp 1738175533
transform 1 0 3680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_30
timestamp 1738175533
transform 1 0 3864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42
timestamp 1738175533
transform 1 0 4968 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1738175533
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1738175533
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1738175533
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1738175533
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1738175533
transform 1 0 5520 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51
timestamp 1738175533
transform 1 0 5796 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1738175533
transform 1 0 6348 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_51
timestamp 1738175533
transform 1 0 5796 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71
timestamp 1738175533
transform 1 0 7636 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_59
timestamp 1738175533
transform 1 0 6532 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_58
timestamp 1738175533
transform 1 0 6440 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_70
timestamp 1738175533
transform 1 0 7544 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1738175533
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output26
timestamp 1738175533
transform -1 0 8648 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77
timestamp 1738175533
transform 1 0 8188 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_82
timestamp 1738175533
transform 1 0 8648 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86
timestamp 1738175533
transform 1 0 9016 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_88
timestamp 1738175533
transform 1 0 9200 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_82
timestamp 1738175533
transform 1 0 8648 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_94
timestamp 1738175533
transform 1 0 9752 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1738175533
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1738175533
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output39
timestamp 1738175533
transform -1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100
timestamp 1738175533
transform 1 0 10304 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1738175533
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_117
timestamp 1738175533
transform 1 0 11868 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_106
timestamp 1738175533
transform 1 0 10856 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_115
timestamp 1738175533
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1738175533
transform -1 0 14076 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_129
timestamp 1738175533
transform 1 0 12972 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_137
timestamp 1738175533
transform 1 0 13708 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1738175533
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_127
timestamp 1738175533
transform 1 0 12788 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_139
timestamp 1738175533
transform 1 0 13892 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1738175533
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output36
timestamp 1738175533
transform 1 0 16376 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_146
timestamp 1738175533
transform 1 0 14536 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_158
timestamp 1738175533
transform 1 0 15640 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_151
timestamp 1738175533
transform 1 0 14996 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_163
timestamp 1738175533
transform 1 0 16100 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1327_
timestamp 1738175533
transform 1 0 17296 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1738175533
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1738175533
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_170
timestamp 1738175533
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1738175533
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1738175533
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1320_
timestamp 1738175533
transform -1 0 18676 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1326_
timestamp 1738175533
transform 1 0 17572 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_182
timestamp 1738175533
transform 1 0 17848 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1738175533
transform 1 0 17664 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1631_
timestamp 1738175533
transform 1 0 18032 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output29
timestamp 1738175533
transform 1 0 19044 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1738175533
transform 1 0 18676 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1738175533
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_200
timestamp 1738175533
transform 1 0 19504 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1319_
timestamp 1738175533
transform 1 0 20424 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1738175533
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_204
timestamp 1738175533
transform 1 0 19872 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_210
timestamp 1738175533
transform 1 0 20424 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_208
timestamp 1738175533
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_214
timestamp 1738175533
transform 1 0 20792 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1632_
timestamp 1738175533
transform 1 0 20516 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _1318_
timestamp 1738175533
transform -1 0 21436 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_221
timestamp 1738175533
transform 1 0 21436 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1738175533
transform 1 0 22448 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1738175533
transform 1 0 22080 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output30
timestamp 1738175533
transform -1 0 23276 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_227
timestamp 1738175533
transform 1 0 21988 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_231
timestamp 1738175533
transform 1 0 22356 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1738175533
transform 1 0 22540 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_227
timestamp 1738175533
transform 1 0 21988 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_229
timestamp 1738175533
transform 1 0 22172 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1738175533
transform 1 0 25116 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_241
timestamp 1738175533
transform 1 0 23276 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1738175533
transform 1 0 24380 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1738175533
transform 1 0 25208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_241
timestamp 1738175533
transform 1 0 23276 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_253
timestamp 1738175533
transform 1 0 24380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1738175533
transform 1 0 27324 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output41
timestamp 1738175533
transform -1 0 25944 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_270
timestamp 1738175533
transform 1 0 25944 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_282
timestamp 1738175533
transform 1 0 27048 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_265
timestamp 1738175533
transform 1 0 25484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_277
timestamp 1738175533
transform 1 0 26588 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_286
timestamp 1738175533
transform 1 0 27416 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _1707_
timestamp 1738175533
transform 1 0 28428 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1738175533
transform 1 0 27784 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output27
timestamp 1738175533
transform -1 0 28612 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_291
timestamp 1738175533
transform 1 0 27876 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_299
timestamp 1738175533
transform 1 0 28612 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_294
timestamp 1738175533
transform 1 0 28152 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1188_
timestamp 1738175533
transform 1 0 30636 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1738175533
transform 1 0 30452 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output33
timestamp 1738175533
transform -1 0 31280 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output37
timestamp 1738175533
transform 1 0 31648 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_311
timestamp 1738175533
transform 1 0 29716 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_320
timestamp 1738175533
transform 1 0 30544 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_328
timestamp 1738175533
transform 1 0 31280 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_317
timestamp 1738175533
transform 1 0 30268 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_324
timestamp 1738175533
transform 1 0 30912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1738175533
transform 1 0 32568 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output35
timestamp 1738175533
transform 1 0 32384 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_336
timestamp 1738175533
transform 1 0 32016 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_344
timestamp 1738175533
transform 1 0 32752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_336
timestamp 1738175533
transform 1 0 32016 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1738175533
transform 1 0 33120 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_349
timestamp 1738175533
transform 1 0 33212 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_357
timestamp 1738175533
transform 1 0 33948 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_355
timestamp 1738175533
transform 1 0 33764 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_343
timestamp 1738175533
transform 1 0 32660 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1738175533
transform -1 0 34316 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1738175533
transform -1 0 34316 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1738175533
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1738175533
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1738175533
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1237_
timestamp 1738175533
transform 1 0 4232 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1738175533
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1738175533
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_30
timestamp 1738175533
transform 1 0 3864 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_43
timestamp 1738175533
transform 1 0 5060 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_47
timestamp 1738175533
transform 1 0 5428 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _1687_
timestamp 1738175533
transform -1 0 7452 0 -1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_2_69
timestamp 1738175533
transform 1 0 7452 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1738175533
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_81
timestamp 1738175533
transform 1 0 8556 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1738175533
transform 1 0 8924 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_87
timestamp 1738175533
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_99
timestamp 1738175533
transform 1 0 10212 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_111
timestamp 1738175533
transform 1 0 11316 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1738175533
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1738175533
transform 1 0 12420 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_135
timestamp 1738175533
transform 1 0 13524 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1628_
timestamp 1738175533
transform -1 0 17572 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_2_144
timestamp 1738175533
transform 1 0 14352 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_156
timestamp 1738175533
transform 1 0 15456 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_162
timestamp 1738175533
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _1321_
timestamp 1738175533
transform 1 0 18124 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_179
timestamp 1738175533
transform 1 0 17572 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_189
timestamp 1738175533
transform 1 0 18492 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1313_
timestamp 1738175533
transform -1 0 21068 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1738175533
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1738175533
transform 1 0 19228 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_201
timestamp 1738175533
transform 1 0 19596 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1738175533
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_217
timestamp 1738175533
transform 1 0 21068 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_229
timestamp 1738175533
transform 1 0 22172 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1738175533
transform 1 0 24748 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_241
timestamp 1738175533
transform 1 0 23276 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_253
timestamp 1738175533
transform 1 0 24380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_258
timestamp 1738175533
transform 1 0 24840 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _1706_
timestamp 1738175533
transform 1 0 26496 0 -1 3808
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_6  FILLER_2_270
timestamp 1738175533
transform 1 0 25944 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1192_
timestamp 1738175533
transform 1 0 29256 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_299
timestamp 1738175533
transform 1 0 28612 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_305
timestamp 1738175533
transform 1 0 29164 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _1191_
timestamp 1738175533
transform -1 0 30820 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _1708_
timestamp 1738175533
transform 1 0 31556 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1738175533
transform 1 0 29992 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_310
timestamp 1738175533
transform 1 0 29624 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_315
timestamp 1738175533
transform 1 0 30084 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_323
timestamp 1738175533
transform 1 0 30820 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_351
timestamp 1738175533
transform 1 0 33396 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_357
timestamp 1738175533
transform 1 0 33948 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1738175533
transform -1 0 34316 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _1685_
timestamp 1738175533
transform 1 0 1932 0 1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1738175533
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1738175533
transform 1 0 1380 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1236_
timestamp 1738175533
transform -1 0 5980 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_30
timestamp 1738175533
transform 1 0 3864 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_42
timestamp 1738175533
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1738175533
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_53
timestamp 1738175533
transform 1 0 5980 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1738175533
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_70
timestamp 1738175533
transform 1 0 7544 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  _1661_
timestamp 1738175533
transform 1 0 9292 0 1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_3_82
timestamp 1738175533
transform 1 0 8648 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_88
timestamp 1738175533
transform 1 0 9200 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1738175533
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_110
timestamp 1738175533
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_115
timestamp 1738175533
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _1658_
timestamp 1738175533
transform -1 0 14812 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_3_127
timestamp 1738175533
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1738175533
transform 1 0 14812 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_161
timestamp 1738175533
transform 1 0 15916 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1738175533
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1738175533
transform 1 0 16652 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_172
timestamp 1738175533
transform 1 0 16928 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_184
timestamp 1738175533
transform 1 0 18032 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1337_
timestamp 1738175533
transform 1 0 20792 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1629_
timestamp 1738175533
transform 1 0 18860 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_3_192
timestamp 1738175533
transform 1 0 18768 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_209
timestamp 1738175533
transform 1 0 20332 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_213
timestamp 1738175533
transform 1 0 20700 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _1730_
timestamp 1738175533
transform 1 0 22632 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1738175533
transform 1 0 22080 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_217
timestamp 1738175533
transform 1 0 21068 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1738175533
transform 1 0 21804 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_229
timestamp 1738175533
transform 1 0 22172 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_233
timestamp 1738175533
transform 1 0 22540 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_254
timestamp 1738175533
transform 1 0 24472 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1738175533
transform 1 0 27324 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_266
timestamp 1738175533
transform 1 0 25576 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_278
timestamp 1738175533
transform 1 0 26680 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_284
timestamp 1738175533
transform 1 0 27232 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_286
timestamp 1738175533
transform 1 0 27416 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1193_
timestamp 1738175533
transform 1 0 28980 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1194_
timestamp 1738175533
transform -1 0 28612 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_3_299
timestamp 1738175533
transform 1 0 28612 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_309
timestamp 1738175533
transform 1 0 29532 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1132_
timestamp 1738175533
transform 1 0 29992 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1189_
timestamp 1738175533
transform 1 0 31188 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_313
timestamp 1738175533
transform 1 0 29900 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_323
timestamp 1738175533
transform 1 0 30820 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_331
timestamp 1738175533
transform 1 0 31556 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1738175533
transform 1 0 32568 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_339
timestamp 1738175533
transform 1 0 32292 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_343
timestamp 1738175533
transform 1 0 32660 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_355
timestamp 1738175533
transform 1 0 33764 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1738175533
transform -1 0 34316 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1238_
timestamp 1738175533
transform 1 0 2576 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1738175533
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output31
timestamp 1738175533
transform -1 0 2116 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1738175533
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_11
timestamp 1738175533
transform 1 0 2116 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_15
timestamp 1738175533
transform 1 0 2484 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _1686_
timestamp 1738175533
transform 1 0 4232 0 -1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1738175533
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_25
timestamp 1738175533
transform 1 0 3404 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_30
timestamp 1738175533
transform 1 0 3864 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_55
timestamp 1738175533
transform 1 0 6164 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_67
timestamp 1738175533
transform 1 0 7268 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1738175533
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_79
timestamp 1738175533
transform 1 0 8372 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 1738175533
transform 1 0 8924 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_87
timestamp 1738175533
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_99
timestamp 1738175533
transform 1 0 10212 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_111
timestamp 1738175533
transform 1 0 11316 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1738175533
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1738175533
transform 1 0 12420 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_135
timestamp 1738175533
transform 1 0 13524 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _1733_
timestamp 1738175533
transform 1 0 14720 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_4_144
timestamp 1738175533
transform 1 0 14352 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1340_
timestamp 1738175533
transform -1 0 18032 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_168
timestamp 1738175533
transform 1 0 16560 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_180
timestamp 1738175533
transform 1 0 17664 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_184
timestamp 1738175533
transform 1 0 18032 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1324_
timestamp 1738175533
transform -1 0 20240 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1325_
timestamp 1738175533
transform 1 0 18768 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1738175533
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_196
timestamp 1738175533
transform 1 0 19136 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_201
timestamp 1738175533
transform 1 0 19596 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_208
timestamp 1738175533
transform 1 0 20240 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1090_
timestamp 1738175533
transform 1 0 22816 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1624_
timestamp 1738175533
transform 1 0 20976 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_232
timestamp 1738175533
transform 1 0 22448 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1738175533
transform 1 0 24748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_245
timestamp 1738175533
transform 1 0 23644 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_258
timestamp 1738175533
transform 1 0 24840 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _1195_
timestamp 1738175533
transform 1 0 27232 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_270
timestamp 1738175533
transform 1 0 25944 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_282
timestamp 1738175533
transform 1 0 27048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_290
timestamp 1738175533
transform 1 0 27784 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_302
timestamp 1738175533
transform 1 0 28888 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1182_
timestamp 1738175533
transform -1 0 30820 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1190_
timestamp 1738175533
transform -1 0 31556 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1738175533
transform 1 0 29992 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_315
timestamp 1738175533
transform 1 0 30084 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_319
timestamp 1738175533
transform 1 0 30452 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_323
timestamp 1738175533
transform 1 0 30820 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_331
timestamp 1738175533
transform 1 0 31556 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1183_
timestamp 1738175533
transform -1 0 32200 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output43
timestamp 1738175533
transform 1 0 33304 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_338
timestamp 1738175533
transform 1 0 32200 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_354
timestamp 1738175533
transform 1 0 33672 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1738175533
transform -1 0 34316 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _1684_
timestamp 1738175533
transform 1 0 1380 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1738175533
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1235_
timestamp 1738175533
transform -1 0 5980 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_24
timestamp 1738175533
transform 1 0 3312 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_36
timestamp 1738175533
transform 1 0 4416 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1738175533
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_53
timestamp 1738175533
transform 1 0 5980 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_58
timestamp 1738175533
transform 1 0 6440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_70
timestamp 1738175533
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1489_
timestamp 1738175533
transform 1 0 9108 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_82
timestamp 1738175533
transform 1 0 8648 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_86
timestamp 1738175533
transform 1 0 9016 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_93
timestamp 1738175533
transform 1 0 9660 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1485_
timestamp 1738175533
transform 1 0 10028 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1738175533
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_104
timestamp 1738175533
transform 1 0 10672 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_112
timestamp 1738175533
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_115
timestamp 1738175533
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1738175533
transform 1 0 13340 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_127
timestamp 1738175533
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_136
timestamp 1738175533
transform 1 0 13616 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1087_
timestamp 1738175533
transform 1 0 15456 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_148
timestamp 1738175533
transform 1 0 14720 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_165
timestamp 1738175533
transform 1 0 16284 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1623_
timestamp 1738175533
transform 1 0 17296 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1738175533
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_172
timestamp 1738175533
transform 1 0 16928 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1338_
timestamp 1738175533
transform 1 0 20608 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_192
timestamp 1738175533
transform 1 0 18768 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_204
timestamp 1738175533
transform 1 0 19872 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1336_
timestamp 1738175533
transform 1 0 21344 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1339_
timestamp 1738175533
transform -1 0 22816 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1738175533
transform 1 0 22080 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_216
timestamp 1738175533
transform 1 0 20976 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_223
timestamp 1738175533
transform 1 0 21620 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_227
timestamp 1738175533
transform 1 0 21988 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_229
timestamp 1738175533
transform 1 0 22172 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_236
timestamp 1738175533
transform 1 0 22816 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1367_
timestamp 1738175533
transform -1 0 23460 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1383_
timestamp 1738175533
transform -1 0 24380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_243
timestamp 1738175533
transform 1 0 23460 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_249
timestamp 1738175533
transform 1 0 24012 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_253
timestamp 1738175533
transform 1 0 24380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1088_
timestamp 1738175533
transform 1 0 25484 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1738175533
transform 1 0 27324 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_274
timestamp 1738175533
transform 1 0 26312 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_282
timestamp 1738175533
transform 1 0 27048 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_286
timestamp 1738175533
transform 1 0 27416 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_298
timestamp 1738175533
transform 1 0 28520 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _1130_
timestamp 1738175533
transform -1 0 31280 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1181_
timestamp 1738175533
transform -1 0 30452 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1187_
timestamp 1738175533
transform -1 0 32016 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_310
timestamp 1738175533
transform 1 0 29624 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_319
timestamp 1738175533
transform 1 0 30452 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_328
timestamp 1738175533
transform 1 0 31280 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1437_
timestamp 1738175533
transform 1 0 33396 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1738175533
transform 1 0 32568 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_336
timestamp 1738175533
transform 1 0 32016 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_343
timestamp 1738175533
transform 1 0 32660 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_354
timestamp 1738175533
transform 1 0 33672 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1738175533
transform -1 0 34316 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1239_
timestamp 1738175533
transform 1 0 2576 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1738175533
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1738175533
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1738175533
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_15
timestamp 1738175533
transform 1 0 2484 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1738175533
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1738175533
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfstp_1  _1689_
timestamp 1738175533
transform 1 0 3864 0 1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1738175533
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_25
timestamp 1738175533
transform 1 0 3404 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1738175533
transform 1 0 3864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_42
timestamp 1738175533
transform 1 0 4968 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_27
timestamp 1738175533
transform 1 0 3588 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1662_
timestamp 1738175533
transform 1 0 6900 0 1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _1688_
timestamp 1738175533
transform -1 0 7544 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1738175533
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_48
timestamp 1738175533
transform 1 0 5520 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_70
timestamp 1738175533
transform 1 0 7544 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_51
timestamp 1738175533
transform 1 0 5796 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_58
timestamp 1738175533
transform 1 0 6440 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_62
timestamp 1738175533
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _0885_
timestamp 1738175533
transform -1 0 10672 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _1490_
timestamp 1738175533
transform -1 0 8648 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1559_
timestamp 1738175533
transform 1 0 9384 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1738175533
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_76
timestamp 1738175533
transform 1 0 8096 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_82
timestamp 1738175533
transform 1 0 8648 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1738175533
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_86
timestamp 1738175533
transform 1 0 9016 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1484_
timestamp 1738175533
transform 1 0 10856 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_104
timestamp 1738175533
transform 1 0 10672 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_99
timestamp 1738175533
transform 1 0 10212 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_105
timestamp 1738175533
transform 1 0 10764 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1738175533
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_112
timestamp 1738175533
transform 1 0 11408 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_109
timestamp 1738175533
transform 1 0 11132 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp 1738175533
transform 1 0 11500 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_115
timestamp 1738175533
transform 1 0 11684 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _1663_
timestamp 1738175533
transform 1 0 11500 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__nand2_1  _1495_
timestamp 1738175533
transform -1 0 12972 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1578_
timestamp 1738175533
transform 1 0 13340 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1738175533
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_133
timestamp 1738175533
transform 1 0 13340 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1738175533
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_123
timestamp 1738175533
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_129
timestamp 1738175533
transform 1 0 12972 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_142
timestamp 1738175533
transform 1 0 14168 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1353_
timestamp 1738175533
transform -1 0 16100 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1619_
timestamp 1738175533
transform 1 0 14812 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_6_144
timestamp 1738175533
transform 1 0 14352 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_156
timestamp 1738175533
transform 1 0 15456 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_163
timestamp 1738175533
transform 1 0 16100 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_148
timestamp 1738175533
transform 1 0 14720 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_165
timestamp 1738175533
transform 1 0 16284 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1341_
timestamp 1738175533
transform 1 0 17296 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1354_
timestamp 1738175533
transform -1 0 16744 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1738175533
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_170
timestamp 1738175533
transform 1 0 16744 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1738175533
transform -1 0 18308 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_180
timestamp 1738175533
transform 1 0 17664 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_184
timestamp 1738175533
transform 1 0 18032 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1618_
timestamp 1738175533
transform -1 0 19596 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_6_187
timestamp 1738175533
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_172
timestamp 1738175533
transform 1 0 16928 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1357_
timestamp 1738175533
transform 1 0 19964 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1363_
timestamp 1738175533
transform -1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1616_
timestamp 1738175533
transform 1 0 19964 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1738175533
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_199
timestamp 1738175533
transform 1 0 19412 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_201
timestamp 1738175533
transform 1 0 19596 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_208
timestamp 1738175533
transform 1 0 20240 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_201
timestamp 1738175533
transform 1 0 19596 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1368_
timestamp 1738175533
transform -1 0 22908 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1615_
timestamp 1738175533
transform 1 0 22080 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1738175533
transform 1 0 22080 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1738175533
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_227
timestamp 1738175533
transform 1 0 21988 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_221
timestamp 1738175533
transform 1 0 21436 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_227
timestamp 1738175533
transform 1 0 21988 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_229
timestamp 1738175533
transform 1 0 22172 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_237
timestamp 1738175533
transform 1 0 22908 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1356_
timestamp 1738175533
transform -1 0 24196 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1365_
timestamp 1738175533
transform -1 0 23920 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1610_
timestamp 1738175533
transform 1 0 24288 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1738175533
transform 1 0 24748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_244
timestamp 1738175533
transform 1 0 23552 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_251
timestamp 1738175533
transform 1 0 24196 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_258
timestamp 1738175533
transform 1 0 24840 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_262
timestamp 1738175533
transform 1 0 25208 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_248
timestamp 1738175533
transform 1 0 23920 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _1732_
timestamp 1738175533
transform 1 0 25300 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1738175533
transform 1 0 27324 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_283
timestamp 1738175533
transform 1 0 27140 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_268
timestamp 1738175533
transform 1 0 25760 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_280
timestamp 1738175533
transform 1 0 26864 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_284
timestamp 1738175533
transform 1 0 27232 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_286
timestamp 1738175533
transform 1 0 27416 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1178_
timestamp 1738175533
transform -1 0 29532 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1180_
timestamp 1738175533
transform 1 0 27876 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _1710_
timestamp 1738175533
transform 1 0 27508 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_6_307
timestamp 1738175533
transform 1 0 29348 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_290
timestamp 1738175533
transform 1 0 27784 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_297
timestamp 1738175533
transform 1 0 28428 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_309
timestamp 1738175533
transform 1 0 29532 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1164_
timestamp 1738175533
transform -1 0 30452 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1738175533
transform 1 0 29992 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_313
timestamp 1738175533
transform 1 0 29900 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_315
timestamp 1738175533
transform 1 0 30084 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_313
timestamp 1738175533
transform 1 0 29900 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1136_
timestamp 1738175533
transform 1 0 30820 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1163_
timestamp 1738175533
transform 1 0 30820 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_327
timestamp 1738175533
transform 1 0 31188 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_319
timestamp 1738175533
transform 1 0 30452 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_326
timestamp 1738175533
transform 1 0 31096 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1184_
timestamp 1738175533
transform 1 0 31464 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_333
timestamp 1738175533
transform 1 0 31740 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_333
timestamp 1738175533
transform 1 0 31740 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1198_
timestamp 1738175533
transform -1 0 33304 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1709_
timestamp 1738175533
transform 1 0 31832 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1738175533
transform 1 0 32568 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_354
timestamp 1738175533
transform 1 0 33672 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_341
timestamp 1738175533
transform 1 0 32476 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_343
timestamp 1738175533
transform 1 0 32660 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_350
timestamp 1738175533
transform 1 0 33304 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1738175533
transform -1 0 34316 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1738175533
transform -1 0 34316 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _1683_
timestamp 1738175533
transform 1 0 1472 0 -1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1738175533
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1738175533
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1234_
timestamp 1738175533
transform 1 0 4876 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1738175533
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_25
timestamp 1738175533
transform 1 0 3404 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_30
timestamp 1738175533
transform 1 0 3864 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_38
timestamp 1738175533
transform 1 0 4600 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_50
timestamp 1738175533
transform 1 0 5704 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_62
timestamp 1738175533
transform 1 0 6808 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1738175533
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_74
timestamp 1738175533
transform 1 0 7912 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_87
timestamp 1738175533
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1562_
timestamp 1738175533
transform 1 0 10672 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_clk_48
timestamp 1738175533
transform -1 0 12236 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_99
timestamp 1738175533
transform 1 0 10212 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_103
timestamp 1738175533
transform 1 0 10580 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_113
timestamp 1738175533
transform 1 0 11500 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_117
timestamp 1738175533
transform 1 0 11868 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1494_
timestamp 1738175533
transform 1 0 13340 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1498_
timestamp 1738175533
transform -1 0 12972 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1738175533
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_121
timestamp 1738175533
transform 1 0 12236 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_125
timestamp 1738175533
transform 1 0 12604 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_129
timestamp 1738175533
transform 1 0 12972 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_138
timestamp 1738175533
transform 1 0 13800 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_142
timestamp 1738175533
transform 1 0 14168 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _1355_
timestamp 1738175533
transform -1 0 15824 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144
timestamp 1738175533
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_160
timestamp 1738175533
transform 1 0 15824 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 1738175533
transform 1 0 16652 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1347_
timestamp 1738175533
transform -1 0 18124 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_168
timestamp 1738175533
transform 1 0 16560 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_172
timestamp 1738175533
transform 1 0 16928 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_180
timestamp 1738175533
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_185
timestamp 1738175533
transform 1 0 18124 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1358_
timestamp 1738175533
transform -1 0 19136 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1364_
timestamp 1738175533
transform -1 0 20700 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1738175533
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_191
timestamp 1738175533
transform 1 0 18676 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_196
timestamp 1738175533
transform 1 0 19136 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_201
timestamp 1738175533
transform 1 0 19596 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_213
timestamp 1738175533
transform 1 0 20700 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1362_
timestamp 1738175533
transform -1 0 21344 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_clk_48
timestamp 1738175533
transform 1 0 21712 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_220
timestamp 1738175533
transform 1 0 21344 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1738175533
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _1384_
timestamp 1738175533
transform 1 0 23736 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1738175533
transform 1 0 24748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_239
timestamp 1738175533
transform 1 0 23092 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_245
timestamp 1738175533
transform 1 0 23644 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_250
timestamp 1738175533
transform 1 0 24104 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_256
timestamp 1738175533
transform 1 0 24656 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_258
timestamp 1738175533
transform 1 0 24840 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _1712_
timestamp 1738175533
transform 1 0 25576 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_8_286
timestamp 1738175533
transform 1 0 27416 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1168_
timestamp 1738175533
transform 1 0 27784 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1177_
timestamp 1738175533
transform 1 0 29348 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1179_
timestamp 1738175533
transform -1 0 28980 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_293
timestamp 1738175533
transform 1 0 28060 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_299
timestamp 1738175533
transform 1 0 28612 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_303
timestamp 1738175533
transform 1 0 28980 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1738175533
transform 1 0 29992 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_310
timestamp 1738175533
transform 1 0 29624 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_315
timestamp 1738175533
transform 1 0 30084 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_327
timestamp 1738175533
transform 1 0 31188 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_333
timestamp 1738175533
transform 1 0 31740 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _1705_
timestamp 1738175533
transform 1 0 31832 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_8_354
timestamp 1738175533
transform 1 0 33672 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1738175533
transform -1 0 34316 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1240_
timestamp 1738175533
transform 1 0 2576 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1738175533
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1738175533
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_15
timestamp 1738175533
transform 1 0 2484 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1233_
timestamp 1738175533
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_25
timestamp 1738175533
transform 1 0 3404 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_37
timestamp 1738175533
transform 1 0 4508 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_43
timestamp 1738175533
transform 1 0 5060 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1530_
timestamp 1738175533
transform 1 0 7176 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1738175533
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_53
timestamp 1738175533
transform 1 0 5980 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_58
timestamp 1738175533
transform 1 0 6440 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1491_
timestamp 1738175533
transform -1 0 8648 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1492_
timestamp 1738175533
transform 1 0 9016 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1529_
timestamp 1738175533
transform 1 0 9752 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_75
timestamp 1738175533
transform 1 0 8004 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_82
timestamp 1738175533
transform 1 0 8648 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_89
timestamp 1738175533
transform 1 0 9292 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_93
timestamp 1738175533
transform 1 0 9660 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1486_
timestamp 1738175533
transform 1 0 10948 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1531_
timestamp 1738175533
transform 1 0 12052 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1738175533
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_103
timestamp 1738175533
transform 1 0 10580 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_110
timestamp 1738175533
transform 1 0 11224 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_115
timestamp 1738175533
transform 1 0 11684 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1496_
timestamp 1738175533
transform 1 0 13616 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_9_128
timestamp 1738175533
transform 1 0 12880 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_141
timestamp 1738175533
transform 1 0 14076 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1361_
timestamp 1738175533
transform -1 0 15916 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1497_
timestamp 1738175533
transform 1 0 14444 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_148
timestamp 1738175533
transform 1 0 14720 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_156
timestamp 1738175533
transform 1 0 15456 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_161
timestamp 1738175533
transform 1 0 15916 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1621_
timestamp 1738175533
transform 1 0 17296 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1738175533
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1738175533
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_172
timestamp 1738175533
transform 1 0 16928 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1351_
timestamp 1738175533
transform -1 0 19872 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_192
timestamp 1738175533
transform 1 0 18768 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_200
timestamp 1738175533
transform 1 0 19504 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_204
timestamp 1738175533
transform 1 0 19872 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1380_
timestamp 1738175533
transform -1 0 22816 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1381_
timestamp 1738175533
transform 1 0 21344 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1738175533
transform 1 0 22080 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_216
timestamp 1738175533
transform 1 0 20976 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_224
timestamp 1738175533
transform 1 0 21712 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_229
timestamp 1738175533
transform 1 0 22172 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_236
timestamp 1738175533
transform 1 0 22816 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1374_
timestamp 1738175533
transform 1 0 24012 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1386_
timestamp 1738175533
transform -1 0 23460 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_clk_48
timestamp 1738175533
transform -1 0 24932 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_243
timestamp 1738175533
transform 1 0 23460 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_252
timestamp 1738175533
transform 1 0 24288 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_259
timestamp 1738175533
transform 1 0 24932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1738175533
transform 1 0 27324 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_271
timestamp 1738175533
transform 1 0 26036 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_283
timestamp 1738175533
transform 1 0 27140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_286
timestamp 1738175533
transform 1 0 27416 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _1172_
timestamp 1738175533
transform 1 0 28704 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1173_
timestamp 1738175533
transform 1 0 27784 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_296
timestamp 1738175533
transform 1 0 28336 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_305
timestamp 1738175533
transform 1 0 29164 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_4  _1133_
timestamp 1738175533
transform 1 0 30544 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_1  _1170_
timestamp 1738175533
transform -1 0 30084 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_311
timestamp 1738175533
transform 1 0 29716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_315
timestamp 1738175533
transform 1 0 30084 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_319
timestamp 1738175533
transform 1 0 30452 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _1174_
timestamp 1738175533
transform 1 0 33028 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1738175533
transform 1 0 32568 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_334
timestamp 1738175533
transform 1 0 31832 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_343
timestamp 1738175533
transform 1 0 32660 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_352
timestamp 1738175533
transform 1 0 33488 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1738175533
transform -1 0 34316 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _1682_
timestamp 1738175533
transform 1 0 1380 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1738175533
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _1690_
timestamp 1738175533
transform 1 0 4508 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1738175533
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1738175533
transform 1 0 3312 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_28
timestamp 1738175533
transform 1 0 3680 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_30
timestamp 1738175533
transform 1 0 3864 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_36
timestamp 1738175533
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _1493_
timestamp 1738175533
transform 1 0 6992 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_58
timestamp 1738175533
transform 1 0 6440 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_68
timestamp 1738175533
transform 1 0 7360 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1488_
timestamp 1738175533
transform -1 0 10028 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1561_
timestamp 1738175533
transform 1 0 7728 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1738175533
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_81
timestamp 1738175533
transform 1 0 8556 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1738175533
transform 1 0 8924 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_87
timestamp 1738175533
transform 1 0 9108 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1499_
timestamp 1738175533
transform -1 0 12236 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1537_
timestamp 1738175533
transform 1 0 10396 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_97
timestamp 1738175533
transform 1 0 10028 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_110
timestamp 1738175533
transform 1 0 11224 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_116
timestamp 1738175533
transform 1 0 11776 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1567_
timestamp 1738175533
transform 1 0 13064 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1738175533
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_121
timestamp 1738175533
transform 1 0 12236 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_129
timestamp 1738175533
transform 1 0 12972 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_139
timestamp 1738175533
transform 1 0 13892 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1617_
timestamp 1738175533
transform 1 0 14720 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_144
timestamp 1738175533
transform 1 0 14352 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_164
timestamp 1738175533
transform 1 0 16192 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1738175533
transform -1 0 18400 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1348_
timestamp 1738175533
transform 1 0 17388 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1359_
timestamp 1738175533
transform -1 0 16836 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_171
timestamp 1738175533
transform 1 0 16836 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_181
timestamp 1738175533
transform 1 0 17756 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_188
timestamp 1738175533
transform 1 0 18400 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _1346_
timestamp 1738175533
transform -1 0 20700 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1738175533
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_201
timestamp 1738175533
transform 1 0 19596 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_213
timestamp 1738175533
transform 1 0 20700 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1611_
timestamp 1738175533
transform 1 0 21344 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1738175533
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_236
timestamp 1738175533
transform 1 0 22816 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1345_
timestamp 1738175533
transform -1 0 23460 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1375_
timestamp 1738175533
transform 1 0 23828 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1738175533
transform 1 0 24748 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_243
timestamp 1738175533
transform 1 0 23460 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_251
timestamp 1738175533
transform 1 0 24196 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_258
timestamp 1738175533
transform 1 0 24840 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_270
timestamp 1738175533
transform 1 0 25944 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_282
timestamp 1738175533
transform 1 0 27048 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1134_
timestamp 1738175533
transform 1 0 27692 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1165_
timestamp 1738175533
transform 1 0 28612 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1175_
timestamp 1738175533
transform -1 0 29624 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_288
timestamp 1738175533
transform 1 0 27600 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_294
timestamp 1738175533
transform 1 0 28152 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_298
timestamp 1738175533
transform 1 0 28520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_302
timestamp 1738175533
transform 1 0 28888 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _1171_
timestamp 1738175533
transform -1 0 31648 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1738175533
transform 1 0 29992 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_310
timestamp 1738175533
transform 1 0 29624 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_315
timestamp 1738175533
transform 1 0 30084 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_332
timestamp 1738175533
transform 1 0 31648 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1131_
timestamp 1738175533
transform -1 0 32936 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1197_
timestamp 1738175533
transform 1 0 33304 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_336
timestamp 1738175533
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_346
timestamp 1738175533
transform 1 0 32936 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_354
timestamp 1738175533
transform 1 0 33672 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1738175533
transform -1 0 34316 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1242_
timestamp 1738175533
transform 1 0 2760 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1738175533
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1738175533
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_6
timestamp 1738175533
transform 1 0 1656 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1231_
timestamp 1738175533
transform 1 0 4232 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_27
timestamp 1738175533
transform 1 0 3588 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_33
timestamp 1738175533
transform 1 0 4140 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_38
timestamp 1738175533
transform 1 0 4600 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1738175533
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_50
timestamp 1738175533
transform 1 0 5704 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_56
timestamp 1738175533
transform 1 0 6256 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_58
timestamp 1738175533
transform 1 0 6440 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_70
timestamp 1738175533
transform 1 0 7544 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1560_
timestamp 1738175533
transform 1 0 8188 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_clk_48
timestamp 1738175533
transform 1 0 9384 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_76
timestamp 1738175533
transform 1 0 8096 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_86
timestamp 1738175533
transform 1 0 9016 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_93
timestamp 1738175533
transform 1 0 9660 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1538_
timestamp 1738175533
transform 1 0 10028 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1738175533
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_clk_48
timestamp 1738175533
transform 1 0 11224 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_106
timestamp 1738175533
transform 1 0 10856 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1738175533
transform 1 0 11500 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_115
timestamp 1738175533
transform 1 0 11684 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1568_
timestamp 1738175533
transform 1 0 12604 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1738175533
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_134
timestamp 1738175533
transform 1 0 13432 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__or2b_1  _0910_
timestamp 1738175533
transform 1 0 15824 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1360_
timestamp 1738175533
transform 1 0 15180 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_146
timestamp 1738175533
transform 1 0 14536 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_152
timestamp 1738175533
transform 1 0 15088 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_156
timestamp 1738175533
transform 1 0 15456 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_166
timestamp 1738175533
transform 1 0 16376 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0916_
timestamp 1738175533
transform -1 0 18032 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1738175533
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk_48
timestamp 1738175533
transform 1 0 17296 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_170
timestamp 1738175533
transform 1 0 16744 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_172
timestamp 1738175533
transform 1 0 16928 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_179
timestamp 1738175533
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_184
timestamp 1738175533
transform 1 0 18032 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_190
timestamp 1738175533
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1316_
timestamp 1738175533
transform -1 0 20884 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1620_
timestamp 1738175533
transform 1 0 18676 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_207
timestamp 1738175533
transform 1 0 20148 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1328_
timestamp 1738175533
transform -1 0 21620 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1350_
timestamp 1738175533
transform -1 0 22908 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1738175533
transform 1 0 22080 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_215
timestamp 1738175533
transform 1 0 20884 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_223
timestamp 1738175533
transform 1 0 21620 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_227
timestamp 1738175533
transform 1 0 21988 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_229
timestamp 1738175533
transform 1 0 22172 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_237
timestamp 1738175533
transform 1 0 22908 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1613_
timestamp 1738175533
transform -1 0 25208 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_clk_48
timestamp 1738175533
transform -1 0 23552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_244
timestamp 1738175533
transform 1 0 23552 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_262
timestamp 1738175533
transform 1 0 25208 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1738175533
transform 1 0 27324 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_274
timestamp 1738175533
transform 1 0 26312 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_282
timestamp 1738175533
transform 1 0 27048 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_286
timestamp 1738175533
transform 1 0 27416 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1169_
timestamp 1738175533
transform 1 0 28152 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1738175533
transform -1 0 29348 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_297
timestamp 1738175533
transform 1 0 28428 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_303
timestamp 1738175533
transform 1 0 28980 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_307
timestamp 1738175533
transform 1 0 29348 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_2  _1162_
timestamp 1738175533
transform 1 0 31372 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1176_
timestamp 1738175533
transform 1 0 29716 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_319
timestamp 1738175533
transform 1 0 30452 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_327
timestamp 1738175533
transform 1 0 31188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_1  _1200_
timestamp 1738175533
transform 1 0 33028 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1738175533
transform 1 0 32568 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_337
timestamp 1738175533
transform 1 0 32108 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_341
timestamp 1738175533
transform 1 0 32476 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_343
timestamp 1738175533
transform 1 0 32660 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_351
timestamp 1738175533
transform 1 0 33396 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_357
timestamp 1738175533
transform 1 0 33948 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1738175533
transform -1 0 34316 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1241_
timestamp 1738175533
transform 1 0 2576 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1738175533
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1738175533
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_15
timestamp 1738175533
transform 1 0 2484 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_23
timestamp 1738175533
transform 1 0 3220 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfstp_1  _1691_
timestamp 1738175533
transform 1 0 4232 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1738175533
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_30
timestamp 1738175533
transform 1 0 3864 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_55
timestamp 1738175533
transform 1 0 6164 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_67
timestamp 1738175533
transform 1 0 7268 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1475_
timestamp 1738175533
transform -1 0 9752 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1480_
timestamp 1738175533
transform -1 0 8648 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1738175533
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_82
timestamp 1738175533
transform 1 0 8648 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1738175533
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_94
timestamp 1738175533
transform 1 0 9752 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1487_
timestamp 1738175533
transform -1 0 10764 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1505_
timestamp 1738175533
transform -1 0 11592 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_105
timestamp 1738175533
transform 1 0 10764 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_114
timestamp 1738175533
transform 1 0 11592 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1502_
timestamp 1738175533
transform 1 0 12604 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1503_
timestamp 1738175533
transform 1 0 13248 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1738175533
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_122
timestamp 1738175533
transform 1 0 12328 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_128
timestamp 1738175533
transform 1 0 12880 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_137
timestamp 1738175533
transform 1 0 13708 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0911_
timestamp 1738175533
transform -1 0 15916 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0912_
timestamp 1738175533
transform 1 0 16284 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_144
timestamp 1738175533
transform 1 0 14352 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_156
timestamp 1738175533
transform 1 0 15456 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_161
timestamp 1738175533
transform 1 0 15916 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0914_
timestamp 1738175533
transform 1 0 17756 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0917_
timestamp 1738175533
transform 1 0 17112 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_168
timestamp 1738175533
transform 1 0 16560 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_177
timestamp 1738175533
transform 1 0 17388 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_187
timestamp 1738175533
transform 1 0 18308 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1331_
timestamp 1738175533
transform -1 0 20792 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1352_
timestamp 1738175533
transform 1 0 18768 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1738175533
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_191
timestamp 1738175533
transform 1 0 18676 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_196
timestamp 1738175533
transform 1 0 19136 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_201
timestamp 1738175533
transform 1 0 19596 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_209
timestamp 1738175533
transform 1 0 20332 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_214
timestamp 1738175533
transform 1 0 20792 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1366_
timestamp 1738175533
transform 1 0 21344 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1370_
timestamp 1738175533
transform 1 0 22540 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_224
timestamp 1738175533
transform 1 0 21712 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_232
timestamp 1738175533
transform 1 0 22448 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_237
timestamp 1738175533
transform 1 0 22908 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1387_
timestamp 1738175533
transform -1 0 23920 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1738175533
transform 1 0 24748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_243
timestamp 1738175533
transform 1 0 23460 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_248
timestamp 1738175533
transform 1 0 23920 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_256
timestamp 1738175533
transform 1 0 24656 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_258
timestamp 1738175533
transform 1 0 24840 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _1711_
timestamp 1738175533
transform 1 0 25668 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_12_266
timestamp 1738175533
transform 1 0 25576 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1135_
timestamp 1738175533
transform 1 0 29348 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1166_
timestamp 1738175533
transform -1 0 28980 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_287
timestamp 1738175533
transform 1 0 27508 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_295
timestamp 1738175533
transform 1 0 28244 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_303
timestamp 1738175533
transform 1 0 28980 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1143_
timestamp 1738175533
transform -1 0 31188 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_4  _1704_
timestamp 1738175533
transform 1 0 31556 0 -1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1738175533
transform 1 0 29992 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_310
timestamp 1738175533
transform 1 0 29624 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_315
timestamp 1738175533
transform 1 0 30084 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_321
timestamp 1738175533
transform 1 0 30636 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_327
timestamp 1738175533
transform 1 0 31188 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_354
timestamp 1738175533
transform 1 0 33672 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1738175533
transform -1 0 34316 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1243_
timestamp 1738175533
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _1681_
timestamp 1738175533
transform 1 0 1380 0 1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1738175533
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1738175533
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1738175533
transform 1 0 1380 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_11
timestamp 1738175533
transform 1 0 2116 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_23
timestamp 1738175533
transform 1 0 3220 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1225_
timestamp 1738175533
transform -1 0 4048 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1232_
timestamp 1738175533
transform 1 0 5060 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1738175533
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_24
timestamp 1738175533
transform 1 0 3312 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_32
timestamp 1738175533
transform 1 0 4048 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_40
timestamp 1738175533
transform 1 0 4784 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1738175533
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_42
timestamp 1738175533
transform 1 0 4968 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1528_
timestamp 1738175533
transform 1 0 6992 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _1660_
timestamp 1738175533
transform 1 0 6808 0 1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1738175533
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1738175533
transform 1 0 5888 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_56
timestamp 1738175533
transform 1 0 6256 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_58
timestamp 1738175533
transform 1 0 6440 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_54
timestamp 1738175533
transform 1 0 6072 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_62
timestamp 1738175533
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_1  _1483_
timestamp 1738175533
transform 1 0 8188 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_73
timestamp 1738175533
transform 1 0 7820 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_81
timestamp 1738175533
transform 1 0 8556 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1474_
timestamp 1738175533
transform 1 0 9476 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1564_
timestamp 1738175533
transform 1 0 9108 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1738175533
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_83
timestamp 1738175533
transform 1 0 8740 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1738175533
transform 1 0 8924 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_87
timestamp 1738175533
transform 1 0 9108 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_94
timestamp 1738175533
transform 1 0 9752 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1476_
timestamp 1738175533
transform 1 0 10304 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1506_
timestamp 1738175533
transform -1 0 10580 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_96
timestamp 1738175533
transform 1 0 9936 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_103
timestamp 1738175533
transform 1 0 10580 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_98
timestamp 1738175533
transform 1 0 10120 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_103
timestamp 1738175533
transform 1 0 10580 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1504_
timestamp 1738175533
transform -1 0 11224 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1536_
timestamp 1738175533
transform 1 0 10948 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1738175533
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_110
timestamp 1738175533
transform 1 0 11224 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115
timestamp 1738175533
transform 1 0 11684 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1535_
timestamp 1738175533
transform 1 0 12052 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_116
timestamp 1738175533
transform 1 0 11776 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1501_
timestamp 1738175533
transform -1 0 13708 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1593_
timestamp 1738175533
transform 1 0 13248 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1738175533
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_clk_48
timestamp 1738175533
transform 1 0 12696 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_128
timestamp 1738175533
transform 1 0 12880 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_141
timestamp 1738175533
transform 1 0 14076 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_124
timestamp 1738175533
transform 1 0 12512 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_129
timestamp 1738175533
transform 1 0 12972 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_137
timestamp 1738175533
transform 1 0 13708 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1334_
timestamp 1738175533
transform 1 0 15548 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1500_
timestamp 1738175533
transform 1 0 14444 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1625_
timestamp 1738175533
transform -1 0 16192 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_13_148
timestamp 1738175533
transform 1 0 14720 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_156
timestamp 1738175533
transform 1 0 15456 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp 1738175533
transform 1 0 15824 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_144
timestamp 1738175533
transform 1 0 14352 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_164
timestamp 1738175533
transform 1 0 16192 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o2111ai_4  _0913_
timestamp 1738175533
transform 1 0 16560 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_2  _0919_
timestamp 1738175533
transform 1 0 17296 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1738175533
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_168
timestamp 1738175533
transform 1 0 16560 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_172
timestamp 1738175533
transform 1 0 16928 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1738175533
transform 1 0 17756 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_189
timestamp 1738175533
transform 1 0 18492 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1343_
timestamp 1738175533
transform 1 0 19688 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1738175533
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_193
timestamp 1738175533
transform 1 0 18860 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_201
timestamp 1738175533
transform 1 0 19596 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1738175533
transform 1 0 19228 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_201
timestamp 1738175533
transform 1 0 19596 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1315_
timestamp 1738175533
transform 1 0 20608 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1344_
timestamp 1738175533
transform -1 0 20332 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_205
timestamp 1738175533
transform 1 0 19964 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_211
timestamp 1738175533
transform 1 0 20516 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1738175533
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1738175533
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1612_
timestamp 1738175533
transform 1 0 20792 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__o21ai_1  _1378_
timestamp 1738175533
transform -1 0 21620 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1738175533
transform 1 0 20884 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_223
timestamp 1738175533
transform 1 0 21620 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1738175533
transform 1 0 22080 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_227
timestamp 1738175533
transform 1 0 21988 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_229
timestamp 1738175533
transform 1 0 22172 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_230
timestamp 1738175533
transform 1 0 22264 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1349_
timestamp 1738175533
transform 1 0 22540 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_clk_48
timestamp 1738175533
transform -1 0 22908 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_236
timestamp 1738175533
transform 1 0 22816 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_237
timestamp 1738175533
transform 1 0 22908 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1342_
timestamp 1738175533
transform -1 0 23368 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1371_
timestamp 1738175533
transform 1 0 23828 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1385_
timestamp 1738175533
transform -1 0 23920 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_244
timestamp 1738175533
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_248
timestamp 1738175533
transform 1 0 23920 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_242
timestamp 1738175533
transform 1 0 23368 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_246
timestamp 1738175533
transform 1 0 23736 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_250
timestamp 1738175533
transform 1 0 24104 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1738175533
transform 1 0 24748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_254
timestamp 1738175533
transform 1 0 24472 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_256
timestamp 1738175533
transform 1 0 24656 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1609_
timestamp 1738175533
transform 1 0 24564 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_14_258
timestamp 1738175533
transform 1 0 24840 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _1713_
timestamp 1738175533
transform 1 0 26588 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1738175533
transform 1 0 27324 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_271
timestamp 1738175533
transform 1 0 26036 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_283
timestamp 1738175533
transform 1 0 27140 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_286
timestamp 1738175533
transform 1 0 27416 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_270
timestamp 1738175533
transform 1 0 25944 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1738175533
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _1137_
timestamp 1738175533
transform -1 0 30084 0 1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_13_298
timestamp 1738175533
transform 1 0 28520 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_297
timestamp 1738175533
transform 1 0 28428 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_309
timestamp 1738175533
transform 1 0 29532 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1167_
timestamp 1738175533
transform 1 0 30452 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1738175533
transform 1 0 29992 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_315
timestamp 1738175533
transform 1 0 30084 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_319
timestamp 1738175533
transform 1 0 30452 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_313
timestamp 1738175533
transform 1 0 29900 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_315
timestamp 1738175533
transform 1 0 30084 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1151_
timestamp 1738175533
transform 1 0 31556 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_13_333
timestamp 1738175533
transform 1 0 31740 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_327
timestamp 1738175533
transform 1 0 31188 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _1144_
timestamp 1738175533
transform -1 0 31740 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _1196_
timestamp 1738175533
transform 1 0 32384 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_14_336
timestamp 1738175533
transform 1 0 32016 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1150_
timestamp 1738175533
transform 1 0 33028 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1738175533
transform 1 0 32568 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_341
timestamp 1738175533
transform 1 0 32476 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_343
timestamp 1738175533
transform 1 0 32660 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_345
timestamp 1738175533
transform 1 0 32844 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1199_
timestamp 1738175533
transform -1 0 33488 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_351
timestamp 1738175533
transform 1 0 33396 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_352
timestamp 1738175533
transform 1 0 33488 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_357
timestamp 1738175533
transform 1 0 33948 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1738175533
transform -1 0 34316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1738175533
transform -1 0 34316 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1226_
timestamp 1738175533
transform -1 0 3588 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1738175533
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1738175533
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_15
timestamp 1738175533
transform 1 0 2484 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfstp_1  _1692_
timestamp 1738175533
transform 1 0 3956 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1738175533
transform 1 0 3588 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1738175533
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1738175533
transform 1 0 5888 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_56
timestamp 1738175533
transform 1 0 6256 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_58
timestamp 1738175533
transform 1 0 6440 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_70
timestamp 1738175533
transform 1 0 7544 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1392_
timestamp 1738175533
transform 1 0 9660 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1565_
timestamp 1738175533
transform 1 0 8188 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_76
timestamp 1738175533
transform 1 0 8096 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_86
timestamp 1738175533
transform 1 0 9016 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_92
timestamp 1738175533
transform 1 0 9568 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1532_
timestamp 1738175533
transform 1 0 10396 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1738175533
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_clk_48
timestamp 1738175533
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_96
timestamp 1738175533
transform 1 0 9936 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_100
timestamp 1738175533
transform 1 0 10304 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_110
timestamp 1738175533
transform 1 0 11224 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_115
timestamp 1738175533
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_2  _0888_
timestamp 1738175533
transform -1 0 13524 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1509_
timestamp 1738175533
transform -1 0 14444 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_122
timestamp 1738175533
transform 1 0 12328 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_126
timestamp 1738175533
transform 1 0 12696 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_135
timestamp 1738175533
transform 1 0 13524 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0915_
timestamp 1738175533
transform 1 0 16192 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1335_
timestamp 1738175533
transform 1 0 15180 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_145
timestamp 1738175533
transform 1 0 14444 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_157
timestamp 1738175533
transform 1 0 15548 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_163
timestamp 1738175533
transform 1 0 16100 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__o2111ai_4  _0918_
timestamp 1738175533
transform 1 0 17480 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1738175533
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_167
timestamp 1738175533
transform 1 0 16468 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_172
timestamp 1738175533
transform 1 0 16928 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1622_
timestamp 1738175533
transform -1 0 21252 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_199
timestamp 1738175533
transform 1 0 19412 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1614_
timestamp 1738175533
transform -1 0 24472 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1738175533
transform 1 0 22080 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_219
timestamp 1738175533
transform 1 0 21252 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_227
timestamp 1738175533
transform 1 0 21988 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_229
timestamp 1738175533
transform 1 0 22172 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_237
timestamp 1738175533
transform 1 0 22908 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _1731_
timestamp 1738175533
transform 1 0 25116 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_15_254
timestamp 1738175533
transform 1 0 24472 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_260
timestamp 1738175533
transform 1 0 25024 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1738175533
transform 1 0 27324 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_281
timestamp 1738175533
transform 1 0 26956 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_286
timestamp 1738175533
transform 1 0 27416 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__o31ai_1  _1156_
timestamp 1738175533
transform -1 0 29624 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_298
timestamp 1738175533
transform 1 0 28520 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _1153_
timestamp 1738175533
transform -1 0 31188 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1160_
timestamp 1738175533
transform 1 0 31556 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_310
timestamp 1738175533
transform 1 0 29624 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_318
timestamp 1738175533
transform 1 0 30360 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_327
timestamp 1738175533
transform 1 0 31188 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1203_
timestamp 1738175533
transform -1 0 33304 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1738175533
transform 1 0 32568 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_335
timestamp 1738175533
transform 1 0 31924 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_341
timestamp 1738175533
transform 1 0 32476 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_343
timestamp 1738175533
transform 1 0 32660 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_350
timestamp 1738175533
transform 1 0 33304 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1738175533
transform -1 0 34316 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _1680_
timestamp 1738175533
transform 1 0 1380 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1738175533
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1230_
timestamp 1738175533
transform 1 0 4876 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1738175533
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1738175533
transform 1 0 3312 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_28
timestamp 1738175533
transform 1 0 3680 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_30
timestamp 1738175533
transform 1 0 3864 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_38
timestamp 1738175533
transform 1 0 4600 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_50
timestamp 1738175533
transform 1 0 5704 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_62
timestamp 1738175533
transform 1 0 6808 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _1512_
timestamp 1738175533
transform -1 0 9936 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1738175533
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_74
timestamp 1738175533
transform 1 0 7912 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1738175533
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _1664_
timestamp 1738175533
transform 1 0 10396 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_16_96
timestamp 1738175533
transform 1 0 9936 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_100
timestamp 1738175533
transform 1 0 10304 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _0886_
timestamp 1738175533
transform 1 0 12696 0 -1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1738175533
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_122
timestamp 1738175533
transform 1 0 12328 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_139
timestamp 1738175533
transform 1 0 13892 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1332_
timestamp 1738175533
transform 1 0 15640 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1508_
timestamp 1738175533
transform -1 0 15180 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_16_144
timestamp 1738175533
transform 1 0 14352 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_153
timestamp 1738175533
transform 1 0 15180 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_157
timestamp 1738175533
transform 1 0 15548 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_161
timestamp 1738175533
transform 1 0 15916 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0897_
timestamp 1738175533
transform -1 0 18308 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0909_
timestamp 1738175533
transform 1 0 16928 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_16_169
timestamp 1738175533
transform 1 0 16652 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_178
timestamp 1738175533
transform 1 0 17480 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_187
timestamp 1738175533
transform 1 0 18308 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1738175533
transform -1 0 19136 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1317_
timestamp 1738175533
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1738175533
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_196
timestamp 1738175533
transform 1 0 19136 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_201
timestamp 1738175533
transform 1 0 19596 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_209
timestamp 1738175533
transform 1 0 20332 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_214
timestamp 1738175533
transform 1 0 20792 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1376_
timestamp 1738175533
transform 1 0 21712 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1377_
timestamp 1738175533
transform -1 0 22632 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_clk_48
timestamp 1738175533
transform -1 0 23276 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_222
timestamp 1738175533
transform 1 0 21528 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_227
timestamp 1738175533
transform 1 0 21988 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_234
timestamp 1738175533
transform 1 0 22632 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1372_
timestamp 1738175533
transform 1 0 23552 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1738175533
transform 1 0 24748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_241
timestamp 1738175533
transform 1 0 23276 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_248
timestamp 1738175533
transform 1 0 23920 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_256
timestamp 1738175533
transform 1 0 24656 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_258
timestamp 1738175533
transform 1 0 24840 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1089_
timestamp 1738175533
transform 1 0 25668 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1373_
timestamp 1738175533
transform -1 0 27140 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_266
timestamp 1738175533
transform 1 0 25576 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_276
timestamp 1738175533
transform 1 0 26496 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_283
timestamp 1738175533
transform 1 0 27140 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _1714_
timestamp 1738175533
transform 1 0 27508 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_16_307
timestamp 1738175533
transform 1 0 29348 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1145_
timestamp 1738175533
transform 1 0 30452 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1152_
timestamp 1738175533
transform -1 0 31372 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1738175533
transform 1 0 29992 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_313
timestamp 1738175533
transform 1 0 29900 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_315
timestamp 1738175533
transform 1 0 30084 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_322
timestamp 1738175533
transform 1 0 30728 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_329
timestamp 1738175533
transform 1 0 31372 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_333
timestamp 1738175533
transform 1 0 31740 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _1703_
timestamp 1738175533
transform 1 0 31832 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_16_354
timestamp 1738175533
transform 1 0 33672 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1738175533
transform -1 0 34316 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1245_
timestamp 1738175533
transform -1 0 3036 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1738175533
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1738175533
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_15
timestamp 1738175533
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_21
timestamp 1738175533
transform 1 0 3036 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1229_
timestamp 1738175533
transform 1 0 4968 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1244_
timestamp 1738175533
transform 1 0 3404 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_28
timestamp 1738175533
transform 1 0 3680 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_40
timestamp 1738175533
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1666_
timestamp 1738175533
transform 1 0 6808 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1738175533
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_51
timestamp 1738175533
transform 1 0 5796 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_58
timestamp 1738175533
transform 1 0 6440 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1573_
timestamp 1738175533
transform 1 0 9108 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_83
timestamp 1738175533
transform 1 0 8740 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1391_
timestamp 1738175533
transform -1 0 10580 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1513_
timestamp 1738175533
transform -1 0 11224 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1738175533
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_96
timestamp 1738175533
transform 1 0 9936 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1738175533
transform 1 0 10580 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_110
timestamp 1738175533
transform 1 0 11224 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_115
timestamp 1738175533
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1596_
timestamp 1738175533
transform 1 0 12880 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_127
timestamp 1738175533
transform 1 0 12788 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_137
timestamp 1738175533
transform 1 0 13708 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1626_
timestamp 1738175533
transform -1 0 15916 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_17_161
timestamp 1738175533
transform 1 0 15916 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1738175533
transform -1 0 17572 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1738175533
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1738175533
transform 1 0 16652 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_172
timestamp 1738175533
transform 1 0 16928 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_179
timestamp 1738175533
transform 1 0 17572 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1627_
timestamp 1738175533
transform 1 0 18952 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_191
timestamp 1738175533
transform 1 0 18676 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_210
timestamp 1738175533
transform 1 0 20424 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1738175533
transform 1 0 22080 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_222
timestamp 1738175533
transform 1 0 21528 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_229
timestamp 1738175533
transform 1 0 22172 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1369_
timestamp 1738175533
transform -1 0 24472 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  repeater45
timestamp 1738175533
transform 1 0 24932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_241
timestamp 1738175533
transform 1 0 23276 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_249
timestamp 1738175533
transform 1 0 24012 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_254
timestamp 1738175533
transform 1 0 24472 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_258
timestamp 1738175533
transform 1 0 24840 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1106_
timestamp 1738175533
transform -1 0 26680 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1738175533
transform 1 0 27324 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_271
timestamp 1738175533
transform 1 0 26036 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_278
timestamp 1738175533
transform 1 0 26680 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_284
timestamp 1738175533
transform 1 0 27232 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_286
timestamp 1738175533
transform 1 0 27416 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1157_
timestamp 1738175533
transform 1 0 29532 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1161_
timestamp 1738175533
transform 1 0 27968 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_298
timestamp 1738175533
transform 1 0 28520 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_306
timestamp 1738175533
transform 1 0 29256 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _1159_
timestamp 1738175533
transform -1 0 31832 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_17_312
timestamp 1738175533
transform 1 0 29808 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1142_
timestamp 1738175533
transform -1 0 33488 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1738175533
transform 1 0 32568 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_334
timestamp 1738175533
transform 1 0 31832 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_343
timestamp 1738175533
transform 1 0 32660 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_352
timestamp 1738175533
transform 1 0 33488 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1738175533
transform -1 0 34316 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1223_
timestamp 1738175533
transform -1 0 3404 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1738175533
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output42
timestamp 1738175533
transform -1 0 2116 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1738175533
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_11
timestamp 1738175533
transform 1 0 2116 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_17
timestamp 1738175533
transform 1 0 2668 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _1693_
timestamp 1738175533
transform 1 0 4600 0 -1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1738175533
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_25
timestamp 1738175533
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_30
timestamp 1738175533
transform 1 0 3864 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_59
timestamp 1738175533
transform 1 0 6532 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_71
timestamp 1738175533
transform 1 0 7636 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1514_
timestamp 1738175533
transform -1 0 8648 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1600_
timestamp 1738175533
transform 1 0 9476 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1738175533
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_82
timestamp 1738175533
transform 1 0 8648 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_87
timestamp 1738175533
transform 1 0 9108 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_100
timestamp 1738175533
transform 1 0 10304 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_112
timestamp 1738175533
transform 1 0 11408 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1507_
timestamp 1738175533
transform -1 0 13340 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1738175533
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_124
timestamp 1738175533
transform 1 0 12512 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_133
timestamp 1738175533
transform 1 0 13340 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1738175533
transform 1 0 14076 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_1  _1333_
timestamp 1738175533
transform 1 0 15364 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_144
timestamp 1738175533
transform 1 0 14352 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_152
timestamp 1738175533
transform 1 0 15088 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_159
timestamp 1738175533
transform 1 0 15732 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0899_
timestamp 1738175533
transform -1 0 17848 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0903_
timestamp 1738175533
transform -1 0 17020 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_167
timestamp 1738175533
transform 1 0 16468 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_173
timestamp 1738175533
transform 1 0 17020 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_182
timestamp 1738175533
transform 1 0 17848 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_190
timestamp 1738175533
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _1329_
timestamp 1738175533
transform -1 0 20240 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1330_
timestamp 1738175533
transform 1 0 18768 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1738175533
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_196
timestamp 1738175533
transform 1 0 19136 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_201
timestamp 1738175533
transform 1 0 19596 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_208
timestamp 1738175533
transform 1 0 20240 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _1728_
timestamp 1738175533
transform -1 0 23092 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_18_216
timestamp 1738175533
transform 1 0 20976 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1097_
timestamp 1738175533
transform 1 0 23460 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1103_
timestamp 1738175533
transform -1 0 24380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1738175533
transform 1 0 24748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_clk_48
timestamp 1738175533
transform -1 0 25484 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_239
timestamp 1738175533
transform 1 0 23092 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_246
timestamp 1738175533
transform 1 0 23736 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_253
timestamp 1738175533
transform 1 0 24380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_258
timestamp 1738175533
transform 1 0 24840 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _1725_
timestamp 1738175533
transform 1 0 25576 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_18_265
timestamp 1738175533
transform 1 0 25484 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_286
timestamp 1738175533
transform 1 0 27416 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1154_
timestamp 1738175533
transform 1 0 29348 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_298
timestamp 1738175533
transform 1 0 28520 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_306
timestamp 1738175533
transform 1 0 29256 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_2  _1146_
timestamp 1738175533
transform -1 0 31280 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1738175533
transform 1 0 29992 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_310
timestamp 1738175533
transform 1 0 29624 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_315
timestamp 1738175533
transform 1 0 30084 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_328
timestamp 1738175533
transform 1 0 31280 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1204_
timestamp 1738175533
transform 1 0 32108 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output34
timestamp 1738175533
transform 1 0 33304 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_336
timestamp 1738175533
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_341
timestamp 1738175533
transform 1 0 32476 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_349
timestamp 1738175533
transform 1 0 33212 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_354
timestamp 1738175533
transform 1 0 33672 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1738175533
transform -1 0 34316 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1227_
timestamp 1738175533
transform 1 0 2484 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _1695_
timestamp 1738175533
transform 1 0 1380 0 1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1738175533
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1738175533
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1738175533
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1228_
timestamp 1738175533
transform -1 0 5428 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1738175533
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_24
timestamp 1738175533
transform 1 0 3312 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1738175533
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1738175533
transform 1 0 5428 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1738175533
transform 1 0 3312 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_28
timestamp 1738175533
transform 1 0 3680 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_30
timestamp 1738175533
transform 1 0 3864 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_42
timestamp 1738175533
transform 1 0 4968 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1534_
timestamp 1738175533
transform 1 0 7452 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _1674_
timestamp 1738175533
transform 1 0 5980 0 -1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1738175533
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_55
timestamp 1738175533
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_58
timestamp 1738175533
transform 1 0 6440 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_66
timestamp 1738175533
transform 1 0 7176 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_50
timestamp 1738175533
transform 1 0 5704 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1516_
timestamp 1738175533
transform -1 0 8648 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_78
timestamp 1738175533
transform 1 0 8280 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_74
timestamp 1738175533
transform 1 0 7912 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1572_
timestamp 1738175533
transform 1 0 8648 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1738175533
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_91
timestamp 1738175533
transform 1 0 9476 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_82
timestamp 1738175533
transform 1 0 8648 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_87
timestamp 1738175533
transform 1 0 9108 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_clk_48
timestamp 1738175533
transform 1 0 9844 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_95
timestamp 1738175533
transform 1 0 9844 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1665_
timestamp 1738175533
transform 1 0 10028 0 -1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1738175533
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1738175533
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_110
timestamp 1738175533
transform 1 0 11224 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_115
timestamp 1738175533
transform 1 0 11684 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1738175533
transform 1 0 12052 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_118
timestamp 1738175533
transform 1 0 11960 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1533_
timestamp 1738175533
transform 1 0 12328 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1598_
timestamp 1738175533
transform 1 0 12604 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_clk_48
timestamp 1738175533
transform -1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1738175533
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_131
timestamp 1738175533
transform 1 0 13156 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1479_
timestamp 1738175533
transform -1 0 13892 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1521_
timestamp 1738175533
transform -1 0 14168 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1738175533
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_134
timestamp 1738175533
transform 1 0 13432 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_139
timestamp 1738175533
transform 1 0 13892 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_142
timestamp 1738175533
transform 1 0 14168 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _0906_
timestamp 1738175533
transform 1 0 16192 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1794_
timestamp 1738175533
transform 1 0 14720 0 -1 13600
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_8  FILLER_19_154
timestamp 1738175533
transform 1 0 15272 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_162
timestamp 1738175533
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_144
timestamp 1738175533
transform 1 0 14352 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o2111ai_4  _0900_
timestamp 1738175533
transform 1 0 17572 0 1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__o2111ai_4  _0907_
timestamp 1738175533
transform 1 0 17204 0 -1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1738175533
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_167
timestamp 1738175533
transform 1 0 16468 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_172
timestamp 1738175533
transform 1 0 16928 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_178
timestamp 1738175533
transform 1 0 17480 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_171
timestamp 1738175533
transform 1 0 16836 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _1724_
timestamp 1738175533
transform 1 0 20056 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1738175533
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_200
timestamp 1738175533
transform 1 0 19504 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_212
timestamp 1738175533
transform 1 0 20608 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_196
timestamp 1738175533
transform 1 0 19136 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_201
timestamp 1738175533
transform 1 0 19596 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_205
timestamp 1738175533
transform 1 0 19964 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_clk_48
timestamp 1738175533
transform 1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_220
timestamp 1738175533
transform 1 0 21344 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1738175533
transform 1 0 22080 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_226
timestamp 1738175533
transform 1 0 21896 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_229
timestamp 1738175533
transform 1 0 22172 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_226
timestamp 1738175533
transform 1 0 21896 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1098_
timestamp 1738175533
transform -1 0 22908 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1118_
timestamp 1738175533
transform 1 0 22724 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_237
timestamp 1738175533
transform 1 0 22908 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_234
timestamp 1738175533
transform 1 0 22632 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _1104_
timestamp 1738175533
transform 1 0 23828 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _1726_
timestamp 1738175533
transform 1 0 23736 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1738175533
transform 1 0 24748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_245
timestamp 1738175533
transform 1 0 23644 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_239
timestamp 1738175533
transform 1 0 23092 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_251
timestamp 1738175533
transform 1 0 24196 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_258
timestamp 1738175533
transform 1 0 24840 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _1107_
timestamp 1738175533
transform 1 0 25944 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_266
timestamp 1738175533
transform 1 0 25576 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_274
timestamp 1738175533
transform 1 0 26312 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_270
timestamp 1738175533
transform 1 0 25944 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1147_
timestamp 1738175533
transform 1 0 26864 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1738175533
transform 1 0 27324 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_282
timestamp 1738175533
transform 1 0 27048 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_286
timestamp 1738175533
transform 1 0 27416 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_278
timestamp 1738175533
transform 1 0 26680 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_284
timestamp 1738175533
transform 1 0 27232 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _1148_
timestamp 1738175533
transform 1 0 28428 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _1716_
timestamp 1738175533
transform 1 0 27784 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_20_296
timestamp 1738175533
transform 1 0 28336 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_303
timestamp 1738175533
transform 1 0 28980 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1149_
timestamp 1738175533
transform -1 0 30728 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1155_
timestamp 1738175533
transform -1 0 30544 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1738175533
transform 1 0 29992 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_310
timestamp 1738175533
transform 1 0 29624 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_320
timestamp 1738175533
transform 1 0 30544 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_311
timestamp 1738175533
transform 1 0 29716 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_315
timestamp 1738175533
transform 1 0 30084 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1158_
timestamp 1738175533
transform 1 0 30912 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1201_
timestamp 1738175533
transform 1 0 31188 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_322
timestamp 1738175533
transform 1 0 30728 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_326
timestamp 1738175533
transform 1 0 31096 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_330
timestamp 1738175533
transform 1 0 31464 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_329
timestamp 1738175533
transform 1 0 31372 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _1206_
timestamp 1738175533
transform 1 0 33028 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _1702_
timestamp 1738175533
transform 1 0 31832 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1738175533
transform 1 0 32568 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_341
timestamp 1738175533
transform 1 0 32476 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_343
timestamp 1738175533
transform 1 0 32660 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_351
timestamp 1738175533
transform 1 0 33396 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_357
timestamp 1738175533
transform 1 0 33948 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_354
timestamp 1738175533
transform 1 0 33672 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1738175533
transform -1 0 34316 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1738175533
transform -1 0 34316 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1738175533
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1738175533
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1738175533
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfstp_1  _1694_
timestamp 1738175533
transform -1 0 5888 0 1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1738175533
transform 1 0 3588 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1390_
timestamp 1738175533
transform -1 0 7084 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1738175533
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1738175533
transform 1 0 5888 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_56
timestamp 1738175533
transform 1 0 6256 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_58
timestamp 1738175533
transform 1 0 6440 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_65
timestamp 1738175533
transform 1 0 7084 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1515_
timestamp 1738175533
transform -1 0 8372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1571_
timestamp 1738175533
transform 1 0 8740 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_73
timestamp 1738175533
transform 1 0 7820 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_79
timestamp 1738175533
transform 1 0 8372 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_92
timestamp 1738175533
transform 1 0 9568 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_8  _1477_
timestamp 1738175533
transform -1 0 13524 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1738175533
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_104
timestamp 1738175533
transform 1 0 10672 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_112
timestamp 1738175533
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_115
timestamp 1738175533
transform 1 0 11684 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1510_
timestamp 1738175533
transform 1 0 13892 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_21_135
timestamp 1738175533
transform 1 0 13524 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1399_
timestamp 1738175533
transform 1 0 16192 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _1526_
timestamp 1738175533
transform -1 0 15824 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_144
timestamp 1738175533
transform 1 0 14352 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_152
timestamp 1738175533
transform 1 0 15088 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_160
timestamp 1738175533
transform 1 0 15824 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1630_
timestamp 1738175533
transform 1 0 17940 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1738175533
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_167
timestamp 1738175533
transform 1 0 16468 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_172
timestamp 1738175533
transform 1 0 16928 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_180
timestamp 1738175533
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1109_
timestamp 1738175533
transform 1 0 20700 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_199
timestamp 1738175533
transform 1 0 19412 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_211
timestamp 1738175533
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _1108_
timestamp 1738175533
transform -1 0 21712 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1721_
timestamp 1738175533
transform 1 0 22632 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1738175533
transform 1 0 22080 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_217
timestamp 1738175533
transform 1 0 21068 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_224
timestamp 1738175533
transform 1 0 21712 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_229
timestamp 1738175533
transform 1 0 22172 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_233
timestamp 1738175533
transform 1 0 22540 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_254
timestamp 1738175533
transform 1 0 24472 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1309_
timestamp 1738175533
transform -1 0 26772 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1738175533
transform 1 0 27324 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_266
timestamp 1738175533
transform 1 0 25576 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_274
timestamp 1738175533
transform 1 0 26312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_279
timestamp 1738175533
transform 1 0 26772 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_286
timestamp 1738175533
transform 1 0 27416 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _1715_
timestamp 1738175533
transform -1 0 31280 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_21_298
timestamp 1738175533
transform 1 0 28520 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_306
timestamp 1738175533
transform 1 0 29256 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  _1186_
timestamp 1738175533
transform 1 0 31648 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_328
timestamp 1738175533
transform 1 0 31280 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1202_
timestamp 1738175533
transform 1 0 33028 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1738175533
transform 1 0 32568 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_336
timestamp 1738175533
transform 1 0 32016 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_343
timestamp 1738175533
transform 1 0 32660 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_352
timestamp 1738175533
transform 1 0 33488 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1738175533
transform -1 0 34316 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0950_
timestamp 1738175533
transform -1 0 3404 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1738175533
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1738175533
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_15
timestamp 1738175533
transform 1 0 2484 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0945_
timestamp 1738175533
transform -1 0 4692 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0953_
timestamp 1738175533
transform -1 0 5428 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1738175533
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_25
timestamp 1738175533
transform 1 0 3404 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_30
timestamp 1738175533
transform 1 0 3864 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_39
timestamp 1738175533
transform 1 0 4692 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_47
timestamp 1738175533
transform 1 0 5428 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1525_
timestamp 1738175533
transform -1 0 7544 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_59
timestamp 1738175533
transform 1 0 6532 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_70
timestamp 1738175533
transform 1 0 7544 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1738175533
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_82
timestamp 1738175533
transform 1 0 8648 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_87
timestamp 1738175533
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _1511_
timestamp 1738175533
transform -1 0 11592 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1599_
timestamp 1738175533
transform 1 0 11960 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_99
timestamp 1738175533
transform 1 0 10212 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_107
timestamp 1738175533
transform 1 0 10948 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_114
timestamp 1738175533
transform 1 0 11592 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1478_
timestamp 1738175533
transform 1 0 13156 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1738175533
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_127
timestamp 1738175533
transform 1 0 12788 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_136
timestamp 1738175533
transform 1 0 13616 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_142
timestamp 1738175533
transform 1 0 14168 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1248_
timestamp 1738175533
transform 1 0 15916 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1527_
timestamp 1738175533
transform 1 0 14996 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_144
timestamp 1738175533
transform 1 0 14352 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_150
timestamp 1738175533
transform 1 0 14904 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_157
timestamp 1738175533
transform 1 0 15548 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_164
timestamp 1738175533
transform 1 0 16192 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _0908_
timestamp 1738175533
transform -1 0 17020 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1323_
timestamp 1738175533
transform 1 0 18032 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_173
timestamp 1738175533
transform 1 0 17020 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_181
timestamp 1738175533
transform 1 0 17756 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_188
timestamp 1738175533
transform 1 0 18400 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1322_
timestamp 1738175533
transform -1 0 19044 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1723_
timestamp 1738175533
transform 1 0 19964 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1738175533
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_195
timestamp 1738175533
transform 1 0 19044 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_199
timestamp 1738175533
transform 1 0 19412 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_201
timestamp 1738175533
transform 1 0 19596 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1096_
timestamp 1738175533
transform 1 0 22908 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1111_
timestamp 1738175533
transform 1 0 22172 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_225
timestamp 1738175533
transform 1 0 21804 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_232
timestamp 1738175533
transform 1 0 22448 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_236
timestamp 1738175533
transform 1 0 22816 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1117_
timestamp 1738175533
transform -1 0 23920 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1738175533
transform 1 0 24748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_241
timestamp 1738175533
transform 1 0 23276 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_248
timestamp 1738175533
transform 1 0 23920 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_256
timestamp 1738175533
transform 1 0 24656 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_258
timestamp 1738175533
transform 1 0 24840 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_262
timestamp 1738175533
transform 1 0 25208 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1307_
timestamp 1738175533
transform -1 0 25576 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1310_
timestamp 1738175533
transform 1 0 25944 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1635_
timestamp 1738175533
transform 1 0 26680 0 -1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_22_266
timestamp 1738175533
transform 1 0 25576 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_274
timestamp 1738175533
transform 1 0 26312 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_295
timestamp 1738175533
transform 1 0 28244 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_307
timestamp 1738175533
transform 1 0 29348 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1214_
timestamp 1738175533
transform -1 0 31004 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1738175533
transform 1 0 29992 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_313
timestamp 1738175533
transform 1 0 29900 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_315
timestamp 1738175533
transform 1 0 30084 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_321
timestamp 1738175533
transform 1 0 30636 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_325
timestamp 1738175533
transform 1 0 31004 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1205_
timestamp 1738175533
transform -1 0 32476 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_337
timestamp 1738175533
transform 1 0 32108 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_341
timestamp 1738175533
transform 1 0 32476 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_353
timestamp 1738175533
transform 1 0 33580 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_357
timestamp 1738175533
transform 1 0 33948 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1738175533
transform -1 0 34316 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1770_
timestamp 1738175533
transform 1 0 1380 0 1 14688
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1738175533
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_2  _0951_
timestamp 1738175533
transform 1 0 3864 0 1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _0952_
timestamp 1738175533
transform -1 0 5796 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_23_26
timestamp 1738175533
transform 1 0 3496 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_40
timestamp 1738175533
transform 1 0 4784 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_8  _0805_
timestamp 1738175533
transform 1 0 7176 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1738175533
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_51
timestamp 1738175533
transform 1 0 5796 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_58
timestamp 1738175533
transform 1 0 6440 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _1775_
timestamp 1738175533
transform -1 0 10856 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_23_82
timestamp 1738175533
transform 1 0 8648 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1482_
timestamp 1738175533
transform -1 0 12420 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1738175533
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_106
timestamp 1738175533
transform 1 0 10856 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_115
timestamp 1738175533
transform 1 0 11684 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1400_
timestamp 1738175533
transform -1 0 14628 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _1401_
timestamp 1738175533
transform 1 0 13064 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_123
timestamp 1738175533
transform 1 0 12420 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_129
timestamp 1738175533
transform 1 0 12972 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1738175533
transform 1 0 13800 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0905_
timestamp 1738175533
transform 1 0 15456 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_23_147
timestamp 1738175533
transform 1 0 14628 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_155
timestamp 1738175533
transform 1 0 15364 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_161
timestamp 1738175533
transform 1 0 15916 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1679_
timestamp 1738175533
transform 1 0 17296 0 1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1738175533
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1738175533
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_172
timestamp 1738175533
transform 1 0 16928 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1112_
timestamp 1738175533
transform 1 0 20608 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_197
timestamp 1738175533
transform 1 0 19228 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_209
timestamp 1738175533
transform 1 0 20332 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1379_
timestamp 1738175533
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1738175533
transform 1 0 22080 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_216
timestamp 1738175533
transform 1 0 20976 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_223
timestamp 1738175533
transform 1 0 21620 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_227
timestamp 1738175533
transform 1 0 21988 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_229
timestamp 1738175533
transform 1 0 22172 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1636_
timestamp 1738175533
transform 1 0 24196 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_23_241
timestamp 1738175533
transform 1 0 23276 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_249
timestamp 1738175533
transform 1 0 24012 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_1  _1305_
timestamp 1738175533
transform 1 0 26496 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1738175533
transform 1 0 27324 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_267
timestamp 1738175533
transform 1 0 25668 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_275
timestamp 1738175533
transform 1 0 26404 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_280
timestamp 1738175533
transform 1 0 26864 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_284
timestamp 1738175533
transform 1 0 27232 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_286
timestamp 1738175533
transform 1 0 27416 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _1698_
timestamp 1738175533
transform 1 0 28980 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_23_298
timestamp 1738175533
transform 1 0 28520 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_302
timestamp 1738175533
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1185_
timestamp 1738175533
transform 1 0 31188 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_323
timestamp 1738175533
transform 1 0 30820 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_330
timestamp 1738175533
transform 1 0 31464 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1209_
timestamp 1738175533
transform 1 0 31832 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1738175533
transform 1 0 32568 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_338
timestamp 1738175533
transform 1 0 32200 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_343
timestamp 1738175533
transform 1 0 32660 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_355
timestamp 1738175533
transform 1 0 33764 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1738175533
transform -1 0 34316 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0949_
timestamp 1738175533
transform 1 0 2852 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1738175533
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1738175533
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_15
timestamp 1738175533
transform 1 0 2484 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _1769_
timestamp 1738175533
transform -1 0 6716 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1738175533
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_25
timestamp 1738175533
transform 1 0 3404 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_30
timestamp 1738175533
transform 1 0 3864 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_38
timestamp 1738175533
transform 1 0 4600 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1524_
timestamp 1738175533
transform -1 0 7912 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_24_61
timestamp 1738175533
transform 1 0 6716 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0947_
timestamp 1738175533
transform -1 0 8648 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1738175533
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_8  repeater46
timestamp 1738175533
transform -1 0 10488 0 -1 15776
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_24_74
timestamp 1738175533
transform 1 0 7912 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_82
timestamp 1738175533
transform 1 0 8648 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_87
timestamp 1738175533
transform 1 0 9108 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0921_
timestamp 1738175533
transform 1 0 10856 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1738175533
transform 1 0 10488 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_113
timestamp 1738175533
transform 1 0 11500 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0889_
timestamp 1738175533
transform -1 0 13708 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0920_
timestamp 1738175533
transform 1 0 12328 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1738175533
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_121
timestamp 1738175533
transform 1 0 12236 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_129
timestamp 1738175533
transform 1 0 12972 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_137
timestamp 1738175533
transform 1 0 13708 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1086_
timestamp 1738175533
transform 1 0 16192 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1247_
timestamp 1738175533
transform -1 0 15824 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_144
timestamp 1738175533
transform 1 0 14352 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_152
timestamp 1738175533
transform 1 0 15088 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_160
timestamp 1738175533
transform 1 0 15824 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1249_
timestamp 1738175533
transform -1 0 17664 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_168
timestamp 1738175533
transform 1 0 16560 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_180
timestamp 1738175533
transform 1 0 17664 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1738175533
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_192
timestamp 1738175533
transform 1 0 18768 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_201
timestamp 1738175533
transform 1 0 19596 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_213
timestamp 1738175533
transform 1 0 20700 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _1722_
timestamp 1738175533
transform 1 0 21712 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_24_221
timestamp 1738175533
transform 1 0 21436 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1308_
timestamp 1738175533
transform -1 0 25576 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1382_
timestamp 1738175533
transform 1 0 23920 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1738175533
transform 1 0 24748 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_244
timestamp 1738175533
transform 1 0 23552 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_251
timestamp 1738175533
transform 1 0 24196 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_258
timestamp 1738175533
transform 1 0 24840 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1105_
timestamp 1738175533
transform -1 0 26220 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1304_
timestamp 1738175533
transform -1 0 27048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_266
timestamp 1738175533
transform 1 0 25576 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_273
timestamp 1738175533
transform 1 0 26220 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_282
timestamp 1738175533
transform 1 0 27048 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1638_
timestamp 1738175533
transform 1 0 27600 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_304
timestamp 1738175533
transform 1 0 29072 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1141_
timestamp 1738175533
transform -1 0 31464 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1738175533
transform 1 0 29992 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_312
timestamp 1738175533
transform 1 0 29808 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_315
timestamp 1738175533
transform 1 0 30084 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_323
timestamp 1738175533
transform 1 0 30820 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_330
timestamp 1738175533
transform 1 0 31464 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _1701_
timestamp 1738175533
transform 1 0 31832 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_24_354
timestamp 1738175533
transform 1 0 33672 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1738175533
transform -1 0 34316 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1771_
timestamp 1738175533
transform 1 0 1380 0 1 15776
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1738175533
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_4  _0799_
timestamp 1738175533
transform -1 0 5336 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_26
timestamp 1738175533
transform 1 0 3496 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_46
timestamp 1738175533
transform 1 0 5336 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1675_
timestamp 1738175533
transform 1 0 7268 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1738175533
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_54
timestamp 1738175533
transform 1 0 6072 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_58
timestamp 1738175533
transform 1 0 6440 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_66
timestamp 1738175533
transform 1 0 7176 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _0893_
timestamp 1738175533
transform 1 0 9660 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_25_88
timestamp 1738175533
transform 1 0 9200 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_92
timestamp 1738175533
transform 1 0 9568 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_1  _0892_
timestamp 1738175533
transform -1 0 11224 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1738175533
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_98
timestamp 1738175533
transform 1 0 10120 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_110
timestamp 1738175533
transform 1 0 11224 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_115
timestamp 1738175533
transform 1 0 11684 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1738175533
transform 1 0 12052 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1246_
timestamp 1738175533
transform 1 0 12880 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1251_
timestamp 1738175533
transform -1 0 14260 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1481_
timestamp 1738175533
transform -1 0 12512 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_124
timestamp 1738175533
transform 1 0 12512 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_131
timestamp 1738175533
transform 1 0 13156 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_137
timestamp 1738175533
transform 1 0 13708 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_143
timestamp 1738175533
transform 1 0 14260 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1738175533
transform -1 0 16100 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1085_
timestamp 1738175533
transform 1 0 14996 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_25_156
timestamp 1738175533
transform 1 0 15456 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_163
timestamp 1738175533
transform 1 0 16100 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1738175533
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_172
timestamp 1738175533
transform 1 0 16928 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_184
timestamp 1738175533
transform 1 0 18032 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_190
timestamp 1738175533
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _1123_
timestamp 1738175533
transform -1 0 19044 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _1719_
timestamp 1738175533
transform -1 0 21344 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_25_195
timestamp 1738175533
transform 1 0 19044 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1115_
timestamp 1738175533
transform 1 0 22540 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1738175533
transform 1 0 22080 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_220
timestamp 1738175533
transform 1 0 21344 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_229
timestamp 1738175533
transform 1 0 22172 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_237
timestamp 1738175533
transform 1 0 22908 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1114_
timestamp 1738175533
transform -1 0 23552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_244
timestamp 1738175533
transform 1 0 23552 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_256
timestamp 1738175533
transform 1 0 24656 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_262
timestamp 1738175533
transform 1 0 25208 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1113_
timestamp 1738175533
transform -1 0 26404 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1116_
timestamp 1738175533
transform -1 0 25760 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1738175533
transform 1 0 27324 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_268
timestamp 1738175533
transform 1 0 25760 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_275
timestamp 1738175533
transform 1 0 26404 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_283
timestamp 1738175533
transform 1 0 27140 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_286
timestamp 1738175533
transform 1 0 27416 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1639_
timestamp 1738175533
transform -1 0 29348 0 1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_25_307
timestamp 1738175533
transform 1 0 29348 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1208_
timestamp 1738175533
transform 1 0 31740 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1213_
timestamp 1738175533
transform 1 0 30084 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_323
timestamp 1738175533
transform 1 0 30820 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_331
timestamp 1738175533
transform 1 0 31556 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1139_
timestamp 1738175533
transform -1 0 33672 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1738175533
transform 1 0 32568 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_338
timestamp 1738175533
transform 1 0 32200 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_343
timestamp 1738175533
transform 1 0 32660 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_354
timestamp 1738175533
transform 1 0 33672 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1738175533
transform -1 0 34316 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0948_
timestamp 1738175533
transform -1 0 3404 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1221_
timestamp 1738175533
transform 1 0 2392 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1738175533
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1738175533
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1738175533
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_15
timestamp 1738175533
transform 1 0 2484 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1738175533
transform 1 0 1380 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_11
timestamp 1738175533
transform 1 0 2116 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_19
timestamp 1738175533
transform 1 0 2852 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__or2b_1  _0801_
timestamp 1738175533
transform -1 0 5244 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1738175533
transform -1 0 5704 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1738175533
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_25
timestamp 1738175533
transform 1 0 3404 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_30
timestamp 1738175533
transform 1 0 3864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_42
timestamp 1738175533
transform 1 0 4968 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_46
timestamp 1738175533
transform 1 0 5336 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_31
timestamp 1738175533
transform 1 0 3956 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_45
timestamp 1738175533
transform 1 0 5244 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0800_
timestamp 1738175533
transform 1 0 5612 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1738175533
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_50
timestamp 1738175533
transform 1 0 5704 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_58
timestamp 1738175533
transform 1 0 6440 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1738175533
transform 1 0 5888 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_56
timestamp 1738175533
transform 1 0 6256 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_58
timestamp 1738175533
transform 1 0 6440 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0807_
timestamp 1738175533
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_27_71
timestamp 1738175533
transform 1 0 7636 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1793_
timestamp 1738175533
transform 1 0 6532 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1653_
timestamp 1738175533
transform 1 0 8188 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1738175533
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_75
timestamp 1738175533
transform 1 0 8004 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_83
timestamp 1738175533
transform 1 0 8740 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1738175533
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _1442_
timestamp 1738175533
transform 1 0 10764 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_27_97
timestamp 1738175533
transform 1 0 10028 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0881_
timestamp 1738175533
transform 1 0 11776 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1738175533
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_111
timestamp 1738175533
transform 1 0 11316 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_115
timestamp 1738175533
transform 1 0 11684 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_119
timestamp 1738175533
transform 1 0 12052 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_110
timestamp 1738175533
transform 1 0 11224 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_115
timestamp 1738175533
transform 1 0 11684 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_99
timestamp 1738175533
transform 1 0 10212 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _0875_
timestamp 1738175533
transform 1 0 13432 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0890_
timestamp 1738175533
transform 1 0 12420 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_4  _0891_
timestamp 1738175533
transform 1 0 12420 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1738175533
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_126
timestamp 1738175533
transform 1 0 12696 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_139
timestamp 1738175533
transform 1 0 13892 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0878_
timestamp 1738175533
transform -1 0 14996 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0880_
timestamp 1738175533
transform 1 0 14720 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_26_144
timestamp 1738175533
transform 1 0 14352 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_151
timestamp 1738175533
transform 1 0 14996 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_144
timestamp 1738175533
transform 1 0 14352 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0874_
timestamp 1738175533
transform -1 0 16284 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0882_
timestamp 1738175533
transform -1 0 16008 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_155
timestamp 1738175533
transform 1 0 15364 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1250_
timestamp 1738175533
transform 1 0 16376 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_162
timestamp 1738175533
transform 1 0 16008 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_165
timestamp 1738175533
transform 1 0 16284 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1433_
timestamp 1738175533
transform -1 0 17296 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1720_
timestamp 1738175533
transform -1 0 19320 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1738175533
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_8  repeater47
timestamp 1738175533
transform -1 0 19136 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_169
timestamp 1738175533
transform 1 0 16652 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_176
timestamp 1738175533
transform 1 0 17296 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_172
timestamp 1738175533
transform 1 0 16928 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_176
timestamp 1738175533
transform 1 0 17296 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1122_
timestamp 1738175533
transform 1 0 19688 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1125_
timestamp 1738175533
transform 1 0 20240 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1738175533
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_196
timestamp 1738175533
transform 1 0 19136 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_201
timestamp 1738175533
transform 1 0 19596 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_207
timestamp 1738175533
transform 1 0 20148 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_212
timestamp 1738175533
transform 1 0 20608 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_198
timestamp 1738175533
transform 1 0 19320 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1738175533
transform 1 0 19964 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _1121_
timestamp 1738175533
transform 1 0 21344 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1124_
timestamp 1738175533
transform 1 0 20976 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1738175533
transform 1 0 22080 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_219
timestamp 1738175533
transform 1 0 21252 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_231
timestamp 1738175533
transform 1 0 22356 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_217
timestamp 1738175533
transform 1 0 21068 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_224
timestamp 1738175533
transform 1 0 21712 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_229
timestamp 1738175533
transform 1 0 22172 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_237
timestamp 1738175533
transform 1 0 22908 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1302_
timestamp 1738175533
transform 1 0 25208 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1727_
timestamp 1738175533
transform -1 0 25024 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1738175533
transform 1 0 24748 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_243
timestamp 1738175533
transform 1 0 23460 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_255
timestamp 1738175533
transform 1 0 24564 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_258
timestamp 1738175533
transform 1 0 24840 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_260
timestamp 1738175533
transform 1 0 25024 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1101_
timestamp 1738175533
transform 1 0 25392 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1110_
timestamp 1738175533
transform -1 0 26312 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_26_265
timestamp 1738175533
transform 1 0 25484 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_274
timestamp 1738175533
transform 1 0 26312 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_272
timestamp 1738175533
transform 1 0 26128 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1102_
timestamp 1738175533
transform -1 0 26772 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1303_
timestamp 1738175533
transform 1 0 26680 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1738175533
transform 1 0 27324 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_279
timestamp 1738175533
transform 1 0 26772 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_286
timestamp 1738175533
transform 1 0 27416 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_282
timestamp 1738175533
transform 1 0 27048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _0963_
timestamp 1738175533
transform 1 0 27968 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1699_
timestamp 1738175533
transform 1 0 28796 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_26_294
timestamp 1738175533
transform 1 0 28152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_306
timestamp 1738175533
transform 1 0 29256 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_295
timestamp 1738175533
transform 1 0 28244 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1138_
timestamp 1738175533
transform 1 0 30452 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1211_
timestamp 1738175533
transform -1 0 32108 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1212_
timestamp 1738175533
transform -1 0 31464 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1738175533
transform 1 0 29992 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_315
timestamp 1738175533
transform 1 0 30084 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_324
timestamp 1738175533
transform 1 0 30912 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_328
timestamp 1738175533
transform 1 0 31280 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_321
timestamp 1738175533
transform 1 0 30636 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_330
timestamp 1738175533
transform 1 0 31464 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1210_
timestamp 1738175533
transform 1 0 31832 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_337
timestamp 1738175533
transform 1 0 32108 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_337
timestamp 1738175533
transform 1 0 32108 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1207_
timestamp 1738175533
transform -1 0 32936 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1738175533
transform 1 0 32568 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_346
timestamp 1738175533
transform 1 0 32936 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_341
timestamp 1738175533
transform 1 0 32476 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_343
timestamp 1738175533
transform 1 0 32660 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1140_
timestamp 1738175533
transform -1 0 33580 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output40
timestamp 1738175533
transform 1 0 33304 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_353
timestamp 1738175533
transform 1 0 33580 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_349
timestamp 1738175533
transform 1 0 33212 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_354
timestamp 1738175533
transform 1 0 33672 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_357
timestamp 1738175533
transform 1 0 33948 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1738175533
transform -1 0 34316 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1738175533
transform -1 0 34316 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1220_
timestamp 1738175533
transform -1 0 2024 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1566_
timestamp 1738175533
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1738175533
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1738175533
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_10
timestamp 1738175533
transform 1 0 2024 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_23
timestamp 1738175533
transform 1 0 3220 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0803_
timestamp 1738175533
transform 1 0 4324 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_4  _0804_
timestamp 1738175533
transform 1 0 4968 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1738175533
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_30
timestamp 1738175533
transform 1 0 3864 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_34
timestamp 1738175533
transform 1 0 4232 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_38
timestamp 1738175533
transform 1 0 4600 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1738175533
transform -1 0 7544 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_63
timestamp 1738175533
transform 1 0 6900 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_70
timestamp 1738175533
transform 1 0 7544 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1738175533
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_82
timestamp 1738175533
transform 1 0 8648 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_87
timestamp 1738175533
transform 1 0 9108 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_95
timestamp 1738175533
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_1  _1650_
timestamp 1738175533
transform 1 0 10028 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_28_118
timestamp 1738175533
transform 1 0 11960 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _0884_
timestamp 1738175533
transform -1 0 13340 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1738175533
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_133
timestamp 1738175533
transform 1 0 13340 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1738175533
transform 1 0 14076 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_2  _1084_
timestamp 1738175533
transform -1 0 15180 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _1654_
timestamp 1738175533
transform 1 0 15548 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_28_144
timestamp 1738175533
transform 1 0 14352 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_153
timestamp 1738175533
transform 1 0 15180 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0873_
timestamp 1738175533
transform 1 0 17756 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_177
timestamp 1738175533
transform 1 0 17388 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_184
timestamp 1738175533
transform 1 0 18032 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _1127_
timestamp 1738175533
transform 1 0 20516 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1738175533
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_196
timestamp 1738175533
transform 1 0 19136 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_201
timestamp 1738175533
transform 1 0 19596 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_209
timestamp 1738175533
transform 1 0 20332 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _1126_
timestamp 1738175533
transform 1 0 21252 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1128_
timestamp 1738175533
transform 1 0 22632 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1129_
timestamp 1738175533
transform 1 0 21896 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1738175533
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_222
timestamp 1738175533
transform 1 0 21528 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_230
timestamp 1738175533
transform 1 0 22264 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_237
timestamp 1738175533
transform 1 0 22908 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1738175533
transform 1 0 24748 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_249
timestamp 1738175533
transform 1 0 24012 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_258
timestamp 1738175533
transform 1 0 24840 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__o22ai_4  _0962_
timestamp 1738175533
transform -1 0 28612 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _0964_
timestamp 1738175533
transform -1 0 26772 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_270
timestamp 1738175533
transform 1 0 25944 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_279
timestamp 1738175533
transform 1 0 26772 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_299
timestamp 1738175533
transform 1 0 28612 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1738175533
transform 1 0 29992 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_311
timestamp 1738175533
transform 1 0 29716 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_315
timestamp 1738175533
transform 1 0 30084 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_327
timestamp 1738175533
transform 1 0 31188 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_333
timestamp 1738175533
transform 1 0 31740 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _1700_
timestamp 1738175533
transform 1 0 31832 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_28_354
timestamp 1738175533
transform 1 0 33672 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1738175533
transform -1 0 34316 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1222_
timestamp 1738175533
transform 1 0 2484 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1738175533
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1738175533
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_22
timestamp 1738175533
transform 1 0 3128 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0946_
timestamp 1738175533
transform 1 0 4692 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1453_
timestamp 1738175533
transform -1 0 4324 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_29_35
timestamp 1738175533
transform 1 0 4324 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_46
timestamp 1738175533
transform 1 0 5336 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_8  _1452_
timestamp 1738175533
transform -1 0 8372 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1738175533
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_54
timestamp 1738175533
transform 1 0 6072 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_58
timestamp 1738175533
transform 1 0 6440 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_62
timestamp 1738175533
transform 1 0 6808 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_1  _1436_
timestamp 1738175533
transform 1 0 8924 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_79
timestamp 1738175533
transform 1 0 8372 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_93
timestamp 1738175533
transform 1 0 9660 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0879_
timestamp 1738175533
transform 1 0 10212 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_4  _1446_
timestamp 1738175533
transform 1 0 12052 0 1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__a21oi_1  _1447_
timestamp 1738175533
transform 1 0 10856 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1738175533
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_102
timestamp 1738175533
transform 1 0 10488 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_110
timestamp 1738175533
transform 1 0 11224 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_115
timestamp 1738175533
transform 1 0 11684 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_140
timestamp 1738175533
transform 1 0 13984 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1738175533
transform -1 0 16468 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_8  _0877_
timestamp 1738175533
transform -1 0 15824 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_160
timestamp 1738175533
transform 1 0 15824 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _1670_
timestamp 1738175533
transform -1 0 19412 0 1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1738175533
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_167
timestamp 1738175533
transform 1 0 16468 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_172
timestamp 1738175533
transform 1 0 16928 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_2  _1718_
timestamp 1738175533
transform -1 0 21712 0 1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_29_199
timestamp 1738175533
transform 1 0 19412 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _1717_
timestamp 1738175533
transform -1 0 24472 0 1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1738175533
transform 1 0 22080 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_224
timestamp 1738175533
transform 1 0 21712 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_229
timestamp 1738175533
transform 1 0 22172 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1640_
timestamp 1738175533
transform 1 0 24840 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_254
timestamp 1738175533
transform 1 0 24472 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1738175533
transform 1 0 27324 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_274
timestamp 1738175533
transform 1 0 26312 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_282
timestamp 1738175533
transform 1 0 27048 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_286
timestamp 1738175533
transform 1 0 27416 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _0966_
timestamp 1738175533
transform -1 0 28980 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_29_303
timestamp 1738175533
transform 1 0 28980 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0828_
timestamp 1738175533
transform 1 0 30360 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_315
timestamp 1738175533
transform 1 0 30084 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_322
timestamp 1738175533
transform 1 0 30728 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1738175533
transform 1 0 32568 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_334
timestamp 1738175533
transform 1 0 31832 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_343
timestamp 1738175533
transform 1 0 32660 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_355
timestamp 1738175533
transform 1 0 33764 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1738175533
transform -1 0 34316 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0797_
timestamp 1738175533
transform -1 0 3404 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0938_
timestamp 1738175533
transform -1 0 2668 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1738175533
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1738175533
transform 1 0 1380 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_11
timestamp 1738175533
transform 1 0 2116 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_17
timestamp 1738175533
transform 1 0 2668 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0927_
timestamp 1738175533
transform -1 0 5152 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1738175533
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_25
timestamp 1738175533
transform 1 0 3404 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_30
timestamp 1738175533
transform 1 0 3864 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_38
timestamp 1738175533
transform 1 0 4600 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_44
timestamp 1738175533
transform 1 0 5152 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0838_
timestamp 1738175533
transform 1 0 5520 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_51
timestamp 1738175533
transform 1 0 5796 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_63
timestamp 1738175533
transform 1 0 6900 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _1422_
timestamp 1738175533
transform -1 0 9936 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1444_
timestamp 1738175533
transform -1 0 8556 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1738175533
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_75
timestamp 1738175533
transform 1 0 8004 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_81
timestamp 1738175533
transform 1 0 8556 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1738175533
transform 1 0 8924 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_87
timestamp 1738175533
transform 1 0 9108 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1443_
timestamp 1738175533
transform 1 0 11500 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1448_
timestamp 1738175533
transform -1 0 10856 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_96
timestamp 1738175533
transform 1 0 9936 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_106
timestamp 1738175533
transform 1 0 10856 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_112
timestamp 1738175533
transform 1 0 11408 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_116
timestamp 1738175533
transform 1 0 11776 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1428_
timestamp 1738175533
transform -1 0 13892 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _1445_
timestamp 1738175533
transform -1 0 12972 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1738175533
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_129
timestamp 1738175533
transform 1 0 12972 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_133
timestamp 1738175533
transform 1 0 13340 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_139
timestamp 1738175533
transform 1 0 13892 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_4  _1427_
timestamp 1738175533
transform 1 0 14904 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_30_144
timestamp 1738175533
transform 1 0 14352 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_166
timestamp 1738175533
transform 1 0 16376 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _1426_
timestamp 1738175533
transform 1 0 18584 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_48
timestamp 1738175533
transform 1 0 16744 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__nand2_2  _1314_
timestamp 1738175533
transform 1 0 19964 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1420_
timestamp 1738175533
transform -1 0 19964 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1738175533
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_197
timestamp 1738175533
transform 1 0 19228 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_210
timestamp 1738175533
transform 1 0 20424 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_222
timestamp 1738175533
transform 1 0 21528 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_234
timestamp 1738175533
transform 1 0 22632 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _1301_
timestamp 1738175533
transform 1 0 25208 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1738175533
transform 1 0 24748 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_246
timestamp 1738175533
transform 1 0 23736 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_254
timestamp 1738175533
transform 1 0 24472 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_258
timestamp 1738175533
transform 1 0 24840 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0961_
timestamp 1738175533
transform -1 0 27232 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1300_
timestamp 1738175533
transform -1 0 26220 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_266
timestamp 1738175533
transform 1 0 25576 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_273
timestamp 1738175533
transform 1 0 26220 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_277
timestamp 1738175533
transform 1 0 26588 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_284
timestamp 1738175533
transform 1 0 27232 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_2  _0965_
timestamp 1738175533
transform 1 0 27876 0 -1 19040
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_30_290
timestamp 1738175533
transform 1 0 27784 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_301
timestamp 1738175533
transform 1 0 28796 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _1763_
timestamp 1738175533
transform 1 0 30452 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1738175533
transform 1 0 29992 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_313
timestamp 1738175533
transform 1 0 29900 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_315
timestamp 1738175533
transform 1 0 30084 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1010_
timestamp 1738175533
transform 1 0 32660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_339
timestamp 1738175533
transform 1 0 32292 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_352
timestamp 1738175533
transform 1 0 33488 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1738175533
transform -1 0 34316 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1773_
timestamp 1738175533
transform 1 0 1380 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1738175533
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_23
timestamp 1738175533
transform 1 0 3220 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0798_
timestamp 1738175533
transform 1 0 3588 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0840_
timestamp 1738175533
transform 1 0 5244 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0940_
timestamp 1738175533
transform 1 0 4508 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_33
timestamp 1738175533
transform 1 0 4140 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 1738175533
transform 1 0 4876 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _1652_
timestamp 1738175533
transform 1 0 6808 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1738175533
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_50
timestamp 1738175533
transform 1 0 5704 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_56
timestamp 1738175533
transform 1 0 6256 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_58
timestamp 1738175533
transform 1 0 6440 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_2  _1429_
timestamp 1738175533
transform -1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_82
timestamp 1738175533
transform 1 0 8648 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1423_
timestamp 1738175533
transform 1 0 10488 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1738175533
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_98
timestamp 1738175533
transform 1 0 10120 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_105
timestamp 1738175533
transform 1 0 10764 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_113
timestamp 1738175533
transform 1 0 11500 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_115
timestamp 1738175533
transform 1 0 11684 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_119
timestamp 1738175533
transform 1 0 12052 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_2  _1255_
timestamp 1738175533
transform 1 0 12144 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1406_
timestamp 1738175533
transform -1 0 13616 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_31_125
timestamp 1738175533
transform 1 0 12604 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_136
timestamp 1738175533
transform 1 0 13616 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1435_
timestamp 1738175533
transform 1 0 15916 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__a41oi_1  _1518_
timestamp 1738175533
transform 1 0 15272 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _1520_
timestamp 1738175533
transform -1 0 15272 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_31_144
timestamp 1738175533
transform 1 0 14352 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _0973_
timestamp 1738175533
transform -1 0 18216 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1738175533
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_167
timestamp 1738175533
transform 1 0 16468 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_172
timestamp 1738175533
transform 1 0 16928 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_186
timestamp 1738175533
transform 1 0 18216 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _1072_
timestamp 1738175533
transform -1 0 21068 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1410_
timestamp 1738175533
transform -1 0 20240 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_31_198
timestamp 1738175533
transform 1 0 19320 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_202
timestamp 1738175533
transform 1 0 19688 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_208
timestamp 1738175533
transform 1 0 20240 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_212
timestamp 1738175533
transform 1 0 20608 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1738175533
transform -1 0 21712 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1071_
timestamp 1738175533
transform 1 0 22540 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1738175533
transform 1 0 22080 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_217
timestamp 1738175533
transform 1 0 21068 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_224
timestamp 1738175533
transform 1 0 21712 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_229
timestamp 1738175533
transform 1 0 22172 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_237
timestamp 1738175533
transform 1 0 22908 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _1736_
timestamp 1738175533
transform 1 0 23276 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_31_261
timestamp 1738175533
transform 1 0 25116 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1065_
timestamp 1738175533
transform 1 0 25484 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1100_
timestamp 1738175533
transform -1 0 26864 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1738175533
transform 1 0 27324 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_269
timestamp 1738175533
transform 1 0 25852 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_275
timestamp 1738175533
transform 1 0 26404 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_280
timestamp 1738175533
transform 1 0 26864 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_284
timestamp 1738175533
transform 1 0 27232 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_286
timestamp 1738175533
transform 1 0 27416 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1634_
timestamp 1738175533
transform -1 0 29900 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_31_294
timestamp 1738175533
transform 1 0 28152 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1011_
timestamp 1738175533
transform 1 0 30544 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_31_313
timestamp 1738175533
transform 1 0 29900 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_319
timestamp 1738175533
transform 1 0 30452 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_329
timestamp 1738175533
transform 1 0 31372 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_1  _0977_
timestamp 1738175533
transform -1 0 33580 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1738175533
transform 1 0 32568 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_341
timestamp 1738175533
transform 1 0 32476 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_343
timestamp 1738175533
transform 1 0 32660 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_353
timestamp 1738175533
transform 1 0 33580 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_357
timestamp 1738175533
transform 1 0 33948 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1738175533
transform -1 0 34316 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0923_
timestamp 1738175533
transform -1 0 3404 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0939_
timestamp 1738175533
transform -1 0 2576 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1738175533
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1738175533
transform 1 0 1380 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_11
timestamp 1738175533
transform 1 0 2116 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_16
timestamp 1738175533
transform 1 0 2576 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0926_
timestamp 1738175533
transform 1 0 4692 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1738175533
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_25
timestamp 1738175533
transform 1 0 3404 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_30
timestamp 1738175533
transform 1 0 3864 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_38
timestamp 1738175533
transform 1 0 4600 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_44
timestamp 1738175533
transform 1 0 5152 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0841_
timestamp 1738175533
transform -1 0 6072 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1738175533
transform 1 0 6716 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_54
timestamp 1738175533
transform 1 0 6072 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_60
timestamp 1738175533
transform 1 0 6624 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_64
timestamp 1738175533
transform 1 0 6992 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__o2111ai_4  _1431_
timestamp 1738175533
transform -1 0 11408 0 -1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1738175533
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_76
timestamp 1738175533
transform 1 0 8096 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_84
timestamp 1738175533
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_87
timestamp 1738175533
transform 1 0 9108 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_112
timestamp 1738175533
transform 1 0 11408 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1254_
timestamp 1738175533
transform 1 0 12972 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1430_
timestamp 1738175533
transform -1 0 12604 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1738175533
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_125
timestamp 1738175533
transform 1 0 12604 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_133
timestamp 1738175533
transform 1 0 13340 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1738175533
transform 1 0 14076 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1425_
timestamp 1738175533
transform -1 0 16100 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1432_
timestamp 1738175533
transform -1 0 15456 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_144
timestamp 1738175533
transform 1 0 14352 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_156
timestamp 1738175533
transform 1 0 15456 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_163
timestamp 1738175533
transform 1 0 16100 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1218_
timestamp 1738175533
transform 1 0 16468 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1434_
timestamp 1738175533
transform 1 0 17572 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_175
timestamp 1738175533
transform 1 0 17204 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_183
timestamp 1738175533
transform 1 0 17940 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _1735_
timestamp 1738175533
transform 1 0 20332 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1738175533
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_195
timestamp 1738175533
transform 1 0 19044 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_199
timestamp 1738175533
transform 1 0 19412 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_201
timestamp 1738175533
transform 1 0 19596 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1070_
timestamp 1738175533
transform 1 0 22632 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_32_229
timestamp 1738175533
transform 1 0 22172 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_233
timestamp 1738175533
transform 1 0 22540 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1738175533
transform -1 0 24380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0968_
timestamp 1738175533
transform -1 0 25668 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1738175533
transform 1 0 24748 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_239
timestamp 1738175533
transform 1 0 23092 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_247
timestamp 1738175533
transform 1 0 23828 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1738175533
transform 1 0 24380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_258
timestamp 1738175533
transform 1 0 24840 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1029_
timestamp 1738175533
transform 1 0 26312 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1099_
timestamp 1738175533
transform 1 0 27048 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_32_267
timestamp 1738175533
transform 1 0 25668 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_273
timestamp 1738175533
transform 1 0 26220 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_278
timestamp 1738175533
transform 1 0 26680 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1311_
timestamp 1738175533
transform -1 0 28980 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_32_287
timestamp 1738175533
transform 1 0 27508 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_293
timestamp 1738175533
transform 1 0 28060 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_303
timestamp 1738175533
transform 1 0 28980 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1738175533
transform 1 0 29992 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_311
timestamp 1738175533
transform 1 0 29716 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_315
timestamp 1738175533
transform 1 0 30084 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_327
timestamp 1738175533
transform 1 0 31188 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_333
timestamp 1738175533
transform 1 0 31740 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _1764_
timestamp 1738175533
transform 1 0 31832 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_32_354
timestamp 1738175533
transform 1 0 33672 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1738175533
transform -1 0 34316 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1738175533
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1738175533
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output28
timestamp 1738175533
transform -1 0 2116 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1738175533
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_11
timestamp 1738175533
transform 1 0 2116 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0937_
timestamp 1738175533
transform 1 0 2944 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0942_
timestamp 1738175533
transform 1 0 2944 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_19
timestamp 1738175533
transform 1 0 2852 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_15
timestamp 1738175533
transform 1 0 2484 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_19
timestamp 1738175533
transform 1 0 2852 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1738175533
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1738175533
transform 1 0 4232 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1738175533
transform 1 0 3864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1738175533
transform 1 0 3772 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_26
timestamp 1738175533
transform 1 0 3496 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_33
timestamp 1738175533
transform 1 0 4140 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp 1738175533
transform 1 0 3312 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_28
timestamp 1738175533
transform 1 0 3680 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_30
timestamp 1738175533
transform 1 0 3864 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1738175533
transform -1 0 5152 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_44
timestamp 1738175533
transform 1 0 5152 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_37
timestamp 1738175533
transform 1 0 4508 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_2  _0928_
timestamp 1738175533
transform 1 0 4876 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1738175533
transform 1 0 6348 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0936_
timestamp 1738175533
transform 1 0 5520 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1738175533
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_51
timestamp 1738175533
transform 1 0 5796 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_58
timestamp 1738175533
transform 1 0 6440 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_53
timestamp 1738175533
transform 1 0 5980 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1450_
timestamp 1738175533
transform 1 0 7176 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_60
timestamp 1738175533
transform 1 0 6624 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_69
timestamp 1738175533
transform 1 0 7452 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _1655_
timestamp 1738175533
transform -1 0 8740 0 1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__a32o_1  _1424_
timestamp 1738175533
transform 1 0 7912 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_73
timestamp 1738175533
transform 1 0 7820 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1738175533
transform 1 0 9016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_83
timestamp 1738175533
transform 1 0 8740 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_82
timestamp 1738175533
transform 1 0 8648 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_87
timestamp 1738175533
transform 1 0 9108 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1282_
timestamp 1738175533
transform 1 0 9568 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1402_
timestamp 1738175533
transform 1 0 9476 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_33_91
timestamp 1738175533
transform 1 0 9476 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_95
timestamp 1738175533
transform 1 0 9844 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o221ai_1  _1403_
timestamp 1738175533
transform 1 0 10488 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1421_
timestamp 1738175533
transform 1 0 10304 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_101
timestamp 1738175533
transform 1 0 10396 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_96
timestamp 1738175533
transform 1 0 9936 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_103
timestamp 1738175533
transform 1 0 10580 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1261_
timestamp 1738175533
transform 1 0 11224 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1738175533
transform 1 0 11592 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_109
timestamp 1738175533
transform 1 0 11132 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_113
timestamp 1738175533
transform 1 0 11500 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_115
timestamp 1738175533
transform 1 0 11684 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_119
timestamp 1738175533
transform 1 0 12052 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_109
timestamp 1738175533
transform 1 0 11132 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_113
timestamp 1738175533
transform 1 0 11500 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_2  _1259_
timestamp 1738175533
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1253_
timestamp 1738175533
transform 1 0 12144 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_123
timestamp 1738175533
transform 1 0 12420 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_131
timestamp 1738175533
transform 1 0 13156 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _1252_
timestamp 1738175533
transform -1 0 14260 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1517_
timestamp 1738175533
transform 1 0 13340 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1738175533
transform 1 0 14260 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_136
timestamp 1738175533
transform 1 0 13616 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1738175533
transform 1 0 14076 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_143
timestamp 1738175533
transform 1 0 14260 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1738175533
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _1216_
timestamp 1738175533
transform 1 0 15732 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _1394_
timestamp 1738175533
transform 1 0 14720 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_1  _1697_
timestamp 1738175533
transform 1 0 16284 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_33_155
timestamp 1738175533
transform 1 0 15364 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_163
timestamp 1738175533
transform 1 0 16100 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_144
timestamp 1738175533
transform 1 0 14352 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_161
timestamp 1738175533
transform 1 0 15916 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1219_
timestamp 1738175533
transform 1 0 18492 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1405_
timestamp 1738175533
transform -1 0 17572 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1696_
timestamp 1738175533
transform 1 0 18032 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1738175533
transform 1 0 16836 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_172
timestamp 1738175533
transform 1 0 16928 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_179
timestamp 1738175533
transform 1 0 17572 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_183
timestamp 1738175533
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_181
timestamp 1738175533
transform 1 0 17756 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_8  _1215_
timestamp 1738175533
transform 1 0 20056 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__or3_1  _1217_
timestamp 1738175533
transform -1 0 20424 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1738175533
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_200
timestamp 1738175533
transform 1 0 19504 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_195
timestamp 1738175533
transform 1 0 19044 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_199
timestamp 1738175533
transform 1 0 19412 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_201
timestamp 1738175533
transform 1 0 19596 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_210
timestamp 1738175533
transform 1 0 20424 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3_4  _1120_
timestamp 1738175533
transform -1 0 24104 0 1 20128
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_1  _1418_
timestamp 1738175533
transform 1 0 22356 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1738175533
transform 1 0 22080 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_222
timestamp 1738175533
transform 1 0 21528 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_229
timestamp 1738175533
transform 1 0 22172 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_235
timestamp 1738175533
transform 1 0 22724 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_222
timestamp 1738175533
transform 1 0 21528 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_230
timestamp 1738175533
transform 1 0 22264 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_234
timestamp 1738175533
transform 1 0 22632 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1066_
timestamp 1738175533
transform 1 0 23276 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_240
timestamp 1738175533
transform 1 0 23184 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_244
timestamp 1738175533
transform 1 0 23552 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1738175533
transform 1 0 23920 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1067_
timestamp 1738175533
transform 1 0 24472 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_250
timestamp 1738175533
transform 1 0 24104 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_251
timestamp 1738175533
transform 1 0 24196 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1738175533
transform 1 0 24748 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_262
timestamp 1738175533
transform 1 0 25208 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_258
timestamp 1738175533
transform 1 0 24840 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0957_
timestamp 1738175533
transform 1 0 25576 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0974_
timestamp 1738175533
transform 1 0 25392 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1024_
timestamp 1738175533
transform 1 0 26404 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1064_
timestamp 1738175533
transform -1 0 26588 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_271
timestamp 1738175533
transform 1 0 26036 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_270
timestamp 1738175533
transform 1 0 25944 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1019_
timestamp 1738175533
transform -1 0 27324 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_279
timestamp 1738175533
transform 1 0 26772 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_277
timestamp 1738175533
transform 1 0 26588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1738175533
transform 1 0 27324 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_286
timestamp 1738175533
transform 1 0 27416 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_285
timestamp 1738175533
transform 1 0 27324 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1312_
timestamp 1738175533
transform 1 0 28060 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1633_
timestamp 1738175533
transform -1 0 29440 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1762_
timestamp 1738175533
transform 1 0 29532 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_33_292
timestamp 1738175533
transform 1 0 27968 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_302
timestamp 1738175533
transform 1 0 28888 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_308
timestamp 1738175533
transform 1 0 29440 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_291
timestamp 1738175533
transform 1 0 27876 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_308
timestamp 1738175533
transform 1 0 29440 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0976_
timestamp 1738175533
transform 1 0 31740 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1012_
timestamp 1738175533
transform 1 0 30452 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1738175533
transform 1 0 29992 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_329
timestamp 1738175533
transform 1 0 31372 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_315
timestamp 1738175533
transform 1 0 30084 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_328
timestamp 1738175533
transform 1 0 31280 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _1761_
timestamp 1738175533
transform 1 0 31832 0 -1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1738175533
transform 1 0 32568 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_338
timestamp 1738175533
transform 1 0 32200 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_343
timestamp 1738175533
transform 1 0 32660 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_355
timestamp 1738175533
transform 1 0 33764 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_354
timestamp 1738175533
transform 1 0 33672 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1738175533
transform -1 0 34316 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1738175533
transform -1 0 34316 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1772_
timestamp 1738175533
transform 1 0 1380 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1738175533
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_23
timestamp 1738175533
transform 1 0 3220 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0941_
timestamp 1738175533
transform -1 0 4140 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1591_
timestamp 1738175533
transform -1 0 5520 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_35_29
timestamp 1738175533
transform 1 0 3772 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_33
timestamp 1738175533
transform 1 0 4140 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1738175533
transform 1 0 6348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_48
timestamp 1738175533
transform 1 0 5520 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_56
timestamp 1738175533
transform 1 0 6256 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_58
timestamp 1738175533
transform 1 0 6440 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_70
timestamp 1738175533
transform 1 0 7544 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__nand3_4  _0871_
timestamp 1738175533
transform -1 0 9016 0 1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__dfrtp_1  _1651_
timestamp 1738175533
transform 1 0 9384 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_35_86
timestamp 1738175533
transform 1 0 9016 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1262_
timestamp 1738175533
transform 1 0 12052 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1738175533
transform 1 0 11592 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_110
timestamp 1738175533
transform 1 0 11224 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_115
timestamp 1738175533
transform 1 0 11684 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o32ai_4  _1396_
timestamp 1738175533
transform 1 0 13800 0 1 21216
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_8  FILLER_35_128
timestamp 1738175533
transform 1 0 12880 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_136
timestamp 1738175533
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_160
timestamp 1738175533
transform 1 0 15824 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0895_
timestamp 1738175533
transform 1 0 17756 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1738175533
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_168
timestamp 1738175533
transform 1 0 16560 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_172
timestamp 1738175533
transform 1 0 16928 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_180
timestamp 1738175533
transform 1 0 17664 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_186
timestamp 1738175533
transform 1 0 18216 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1738175533
transform -1 0 20148 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_198
timestamp 1738175533
transform 1 0 19320 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_207
timestamp 1738175533
transform 1 0 20148 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_1  _1411_
timestamp 1738175533
transform -1 0 21712 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1419_
timestamp 1738175533
transform -1 0 23276 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1738175533
transform 1 0 22080 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_224
timestamp 1738175533
transform 1 0 21712 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_229
timestamp 1738175533
transform 1 0 22172 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1439_
timestamp 1738175533
transform 1 0 24380 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_241
timestamp 1738175533
transform 1 0 23276 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_259
timestamp 1738175533
transform 1 0 24932 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0972_
timestamp 1738175533
transform -1 0 25760 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1738175533
transform 1 0 27324 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_268
timestamp 1738175533
transform 1 0 25760 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_280
timestamp 1738175533
transform 1 0 26864 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_284
timestamp 1738175533
transform 1 0 27232 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_286
timestamp 1738175533
transform 1 0 27416 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1018_
timestamp 1738175533
transform -1 0 28612 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1023_
timestamp 1738175533
transform -1 0 29348 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_299
timestamp 1738175533
transform 1 0 28612 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_307
timestamp 1738175533
transform 1 0 29348 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1009_
timestamp 1738175533
transform 1 0 30360 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1013_
timestamp 1738175533
transform -1 0 32200 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_35_315
timestamp 1738175533
transform 1 0 30084 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_322
timestamp 1738175533
transform 1 0 30728 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_328
timestamp 1738175533
transform 1 0 31280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1738175533
transform 1 0 32568 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1738175533
transform -1 0 33672 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_338
timestamp 1738175533
transform 1 0 32200 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_343
timestamp 1738175533
transform 1 0 32660 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_354
timestamp 1738175533
transform 1 0 33672 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1738175533
transform -1 0 34316 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0944_
timestamp 1738175533
transform -1 0 3036 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1738175533
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1738175533
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_15
timestamp 1738175533
transform 1 0 2484 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_21
timestamp 1738175533
transform 1 0 3036 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0934_
timestamp 1738175533
transform 1 0 4692 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1441_
timestamp 1738175533
transform -1 0 5612 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1738175533
transform 1 0 3772 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_30
timestamp 1738175533
transform 1 0 3864 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_38
timestamp 1738175533
transform 1 0 4600 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_42
timestamp 1738175533
transform 1 0 4968 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _0867_
timestamp 1738175533
transform -1 0 7544 0 -1 22304
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_36_49
timestamp 1738175533
transform 1 0 5612 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_55
timestamp 1738175533
transform 1 0 6164 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_70
timestamp 1738175533
transform 1 0 7544 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1738175533
transform 1 0 9016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_82
timestamp 1738175533
transform 1 0 8648 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_87
timestamp 1738175533
transform 1 0 9108 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0872_
timestamp 1738175533
transform -1 0 11224 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _1260_
timestamp 1738175533
transform -1 0 12604 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_36_99
timestamp 1738175533
transform 1 0 10212 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_105
timestamp 1738175533
transform 1 0 10764 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_110
timestamp 1738175533
transform 1 0 11224 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1519_
timestamp 1738175533
transform 1 0 13340 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1738175533
transform 1 0 14260 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_125
timestamp 1738175533
transform 1 0 12604 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_137
timestamp 1738175533
transform 1 0 13708 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1451_
timestamp 1738175533
transform 1 0 16284 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_36_144
timestamp 1738175533
transform 1 0 14352 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_156
timestamp 1738175533
transform 1 0 15456 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_164
timestamp 1738175533
transform 1 0 16192 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_170
timestamp 1738175533
transform 1 0 16744 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_182
timestamp 1738175533
transform 1 0 17848 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _1668_
timestamp 1738175533
transform 1 0 20148 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1738175533
transform 1 0 19504 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_194
timestamp 1738175533
transform 1 0 18952 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_201
timestamp 1738175533
transform 1 0 19596 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_4  _0980_
timestamp 1738175533
transform -1 0 23828 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_227
timestamp 1738175533
transform 1 0 21988 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1738175533
transform 1 0 24748 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_247
timestamp 1738175533
transform 1 0 23828 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_255
timestamp 1738175533
transform 1 0 24564 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_258
timestamp 1738175533
transform 1 0 24840 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__o2111ai_4  _0979_
timestamp 1738175533
transform -1 0 27876 0 -1 22304
box -38 -48 1970 592
use sky130_fd_sc_hd__nand3_4  _1063_
timestamp 1738175533
transform 1 0 28244 0 -1 22304
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_36_291
timestamp 1738175533
transform 1 0 27876 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_309
timestamp 1738175533
transform 1 0 29532 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0975_
timestamp 1738175533
transform 1 0 30636 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_4  _0978_
timestamp 1738175533
transform -1 0 32752 0 -1 22304
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1738175533
transform 1 0 29992 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_313
timestamp 1738175533
transform 1 0 29900 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_315
timestamp 1738175533
transform 1 0 30084 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_326
timestamp 1738175533
transform 1 0 31096 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_344
timestamp 1738175533
transform 1 0 32752 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_356
timestamp 1738175533
transform 1 0 33856 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1738175533
transform -1 0 34316 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0943_
timestamp 1738175533
transform -1 0 2944 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1738175533
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1738175533
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_15
timestamp 1738175533
transform 1 0 2484 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_20
timestamp 1738175533
transform 1 0 2944 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0831_
timestamp 1738175533
transform -1 0 3588 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0935_
timestamp 1738175533
transform 1 0 4140 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_27
timestamp 1738175533
transform 1 0 3588 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_41
timestamp 1738175533
transform 1 0 4876 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_47
timestamp 1738175533
transform 1 0 5428 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _0931_
timestamp 1738175533
transform 1 0 5520 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _1734_
timestamp 1738175533
transform -1 0 8740 0 1 22304
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1738175533
transform 1 0 6348 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_53
timestamp 1738175533
transform 1 0 5980 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_58
timestamp 1738175533
transform 1 0 6440 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1074_
timestamp 1738175533
transform 1 0 9108 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_83
timestamp 1738175533
transform 1 0 8740 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_91
timestamp 1738175533
transform 1 0 9476 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1080_
timestamp 1738175533
transform -1 0 11132 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1258_
timestamp 1738175533
transform 1 0 12052 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1738175533
transform 1 0 11592 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_103
timestamp 1738175533
transform 1 0 10580 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_109
timestamp 1738175533
transform 1 0 11132 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_113
timestamp 1738175533
transform 1 0 11500 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_115
timestamp 1738175533
transform 1 0 11684 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1407_
timestamp 1738175533
transform 1 0 12880 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _1657_
timestamp 1738175533
transform 1 0 14076 0 1 22304
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_37_122
timestamp 1738175533
transform 1 0 12328 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_132
timestamp 1738175533
transform 1 0 13248 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_140
timestamp 1738175533
transform 1 0 13984 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_162
timestamp 1738175533
transform 1 0 16008 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _1768_
timestamp 1738175533
transform -1 0 19136 0 1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1738175533
transform 1 0 16836 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_170
timestamp 1738175533
transform 1 0 16744 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_172
timestamp 1738175533
transform 1 0 16928 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _0998_
timestamp 1738175533
transform -1 0 19964 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_1  _1094_
timestamp 1738175533
transform 1 0 20332 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_37_196
timestamp 1738175533
transform 1 0 19136 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_205
timestamp 1738175533
transform 1 0 19964 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_214
timestamp 1738175533
transform 1 0 20792 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _0994_
timestamp 1738175533
transform -1 0 23000 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1738175533
transform 1 0 22080 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_226
timestamp 1738175533
transform 1 0 21896 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_229
timestamp 1738175533
transform 1 0 22172 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_238
timestamp 1738175533
transform 1 0 23000 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2ai_1  _1440_
timestamp 1738175533
transform 1 0 23368 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_2  _1669_
timestamp 1738175533
transform 1 0 24380 0 1 22304
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_37_249
timestamp 1738175533
transform 1 0 24012 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1738175533
transform 1 0 26680 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1738175533
transform 1 0 27324 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_274
timestamp 1738175533
transform 1 0 26312 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_281
timestamp 1738175533
transform 1 0 26956 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_286
timestamp 1738175533
transform 1 0 27416 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _1758_
timestamp 1738175533
transform 1 0 28244 0 1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_37_294
timestamp 1738175533
transform 1 0 28152 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1015_
timestamp 1738175533
transform 1 0 30820 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_37_315
timestamp 1738175533
transform 1 0 30084 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_332
timestamp 1738175533
transform 1 0 31648 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1738175533
transform 1 0 32568 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_340
timestamp 1738175533
transform 1 0 32384 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_343
timestamp 1738175533
transform 1 0 32660 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_355
timestamp 1738175533
transform 1 0 33764 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1738175533
transform -1 0 34316 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1774_
timestamp 1738175533
transform 1 0 1380 0 -1 23392
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1738175533
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_4  _0932_
timestamp 1738175533
transform -1 0 6348 0 -1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1738175533
transform 1 0 3772 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1738175533
transform 1 0 3312 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_28
timestamp 1738175533
transform 1 0 3680 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_30
timestamp 1738175533
transform 1 0 3864 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_38
timestamp 1738175533
transform 1 0 4600 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_8  _0868_
timestamp 1738175533
transform 1 0 6900 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_38_57
timestamp 1738175533
transform 1 0 6348 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1738175533
transform 1 0 9016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_79
timestamp 1738175533
transform 1 0 8372 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_85
timestamp 1738175533
transform 1 0 8924 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_87
timestamp 1738175533
transform 1 0 9108 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_95
timestamp 1738175533
transform 1 0 9844 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__o31ai_2  _1079_
timestamp 1738175533
transform -1 0 10948 0 -1 23392
box -38 -48 958 592
use sky130_fd_sc_hd__nand3_1  _1266_
timestamp 1738175533
transform 1 0 11868 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_107
timestamp 1738175533
transform 1 0 10948 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_115
timestamp 1738175533
transform 1 0 11684 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _1257_
timestamp 1738175533
transform -1 0 12880 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1738175533
transform 1 0 14260 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_121
timestamp 1738175533
transform 1 0 12236 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_128
timestamp 1738175533
transform 1 0 12880 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_140
timestamp 1738175533
transform 1 0 13984 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1395_
timestamp 1738175533
transform -1 0 14996 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1765_
timestamp 1738175533
transform 1 0 15824 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_144
timestamp 1738175533
transform 1 0 14352 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_151
timestamp 1738175533
transform 1 0 14996 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_159
timestamp 1738175533
transform 1 0 15732 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1002_
timestamp 1738175533
transform 1 0 17664 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_176
timestamp 1738175533
transform 1 0 17296 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_184
timestamp 1738175533
transform 1 0 18032 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0999_
timestamp 1738175533
transform 1 0 18768 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1417_
timestamp 1738175533
transform 1 0 20332 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1738175533
transform 1 0 19504 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_196
timestamp 1738175533
transform 1 0 19136 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_201
timestamp 1738175533
transform 1 0 19596 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_8  repeater48
timestamp 1738175533
transform -1 0 22448 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_216
timestamp 1738175533
transform 1 0 20976 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_232
timestamp 1738175533
transform 1 0 22448 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1119_
timestamp 1738175533
transform -1 0 23828 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1738175533
transform 1 0 24748 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_240
timestamp 1738175533
transform 1 0 23184 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_247
timestamp 1738175533
transform 1 0 23828 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_255
timestamp 1738175533
transform 1 0 24564 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_258
timestamp 1738175533
transform 1 0 24840 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_262
timestamp 1738175533
transform 1 0 25208 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1306_
timestamp 1738175533
transform 1 0 25300 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_38_272
timestamp 1738175533
transform 1 0 26128 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_284
timestamp 1738175533
transform 1 0 27232 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0809_
timestamp 1738175533
transform -1 0 27876 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1017_
timestamp 1738175533
transform 1 0 28336 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_38_291
timestamp 1738175533
transform 1 0 27876 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_295
timestamp 1738175533
transform 1 0 28244 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_305
timestamp 1738175533
transform 1 0 29164 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _1759_
timestamp 1738175533
transform 1 0 30636 0 -1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1738175533
transform 1 0 29992 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_313
timestamp 1738175533
transform 1 0 29900 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_315
timestamp 1738175533
transform 1 0 30084 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1014_
timestamp 1738175533
transform 1 0 32844 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_38_341
timestamp 1738175533
transform 1 0 32476 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_354
timestamp 1738175533
transform 1 0 33672 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1738175533
transform -1 0 34316 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0862_
timestamp 1738175533
transform 1 0 2116 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1738175533
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1738175533
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1738175533
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_6
timestamp 1738175533
transform 1 0 1656 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_10
timestamp 1738175533
transform 1 0 2024 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0832_
timestamp 1738175533
transform 1 0 3220 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1738175533
transform -1 0 2852 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1224_
timestamp 1738175533
transform -1 0 3404 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_39_15
timestamp 1738175533
transform 1 0 2484 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_19
timestamp 1738175533
transform 1 0 2852 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_14
timestamp 1738175533
transform 1 0 2392 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1738175533
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_4  _0929_
timestamp 1738175533
transform 1 0 4416 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__o211ai_4  _0933_
timestamp 1738175533
transform -1 0 5980 0 1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1738175533
transform 1 0 3772 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_27
timestamp 1738175533
transform 1 0 3588 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_35
timestamp 1738175533
transform 1 0 4324 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_25
timestamp 1738175533
transform 1 0 3404 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_30
timestamp 1738175533
transform 1 0 3864 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1738175533
transform 1 0 6164 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1738175533
transform 1 0 6348 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_53
timestamp 1738175533
transform 1 0 5980 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_58
timestamp 1738175533
transform 1 0 6440 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1738175533
transform 1 0 7544 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_49
timestamp 1738175533
transform 1 0 5612 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_58
timestamp 1738175533
transform 1 0 6440 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_70
timestamp 1738175533
transform 1 0 7544 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _0870_
timestamp 1738175533
transform 1 0 8004 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1081_
timestamp 1738175533
transform 1 0 8740 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1083_
timestamp 1738175533
transform -1 0 8372 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_74
timestamp 1738175533
transform 1 0 7912 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_79
timestamp 1738175533
transform 1 0 8372 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_74
timestamp 1738175533
transform 1 0 7912 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_80
timestamp 1738175533
transform 1 0 8464 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1082_
timestamp 1738175533
transform -1 0 10028 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1738175533
transform 1 0 9016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1738175533
transform 1 0 9384 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_87
timestamp 1738175533
transform 1 0 9108 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_93
timestamp 1738175533
transform 1 0 9660 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _1677_
timestamp 1738175533
transform -1 0 11592 0 -1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__nand2_1  _1268_
timestamp 1738175533
transform -1 0 10672 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1738175533
transform 1 0 11592 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_97
timestamp 1738175533
transform 1 0 10028 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_104
timestamp 1738175533
transform 1 0 10672 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_112
timestamp 1738175533
transform 1 0 11408 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_115
timestamp 1738175533
transform 1 0 11684 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_119
timestamp 1738175533
transform 1 0 12052 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_114
timestamp 1738175533
transform 1 0 11592 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1263_
timestamp 1738175533
transform -1 0 12512 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1264_
timestamp 1738175533
transform 1 0 12144 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1265_
timestamp 1738175533
transform 1 0 12880 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1678_
timestamp 1738175533
transform 1 0 13156 0 1 23392
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1738175533
transform 1 0 14260 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_124
timestamp 1738175533
transform 1 0 12512 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_130
timestamp 1738175533
transform 1 0 13064 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_124
timestamp 1738175533
transform 1 0 12512 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_131
timestamp 1738175533
transform 1 0 13156 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2b_1  _1008_
timestamp 1738175533
transform -1 0 16560 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_39_152
timestamp 1738175533
transform 1 0 15088 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_164
timestamp 1738175533
transform 1 0 16192 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_144
timestamp 1738175533
transform 1 0 14352 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_156
timestamp 1738175533
transform 1 0 15456 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_162
timestamp 1738175533
transform 1 0 16008 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _1006_
timestamp 1738175533
transform 1 0 16928 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1738175533
transform 1 0 16836 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_170
timestamp 1738175533
transform 1 0 16744 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_168
timestamp 1738175533
transform 1 0 16560 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1007_
timestamp 1738175533
transform 1 0 17940 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_179
timestamp 1738175533
transform 1 0 17572 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_186
timestamp 1738175533
transform 1 0 18216 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_190
timestamp 1738175533
transform 1 0 18584 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_172
timestamp 1738175533
transform 1 0 16928 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1738175533
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0996_
timestamp 1738175533
transform 1 0 19964 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1003_
timestamp 1738175533
transform -1 0 19136 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1095_
timestamp 1738175533
transform 1 0 19412 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1738175533
transform 1 0 19504 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_196
timestamp 1738175533
transform 1 0 19136 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_203
timestamp 1738175533
transform 1 0 19780 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_196
timestamp 1738175533
transform 1 0 19136 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_201
timestamp 1738175533
transform 1 0 19596 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_209
timestamp 1738175533
transform 1 0 20332 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfstp_1  _1667_
timestamp 1738175533
transform 1 0 20976 0 -1 24480
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1738175533
transform 1 0 22080 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_clk_48
timestamp 1738175533
transform 1 0 22724 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_215
timestamp 1738175533
transform 1 0 20884 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_227
timestamp 1738175533
transform 1 0 21988 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_229
timestamp 1738175533
transform 1 0 22172 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_238
timestamp 1738175533
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_215
timestamp 1738175533
transform 1 0 20884 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_237
timestamp 1738175533
transform 1 0 22908 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1016_
timestamp 1738175533
transform 1 0 24104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1438_
timestamp 1738175533
transform 1 0 23276 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_40_246
timestamp 1738175533
transform 1 0 23736 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1738175533
transform 1 0 24748 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_clk_48
timestamp 1738175533
transform -1 0 25392 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_254
timestamp 1738175533
transform 1 0 24472 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_260
timestamp 1738175533
transform 1 0 25024 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_253
timestamp 1738175533
transform 1 0 24380 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_258
timestamp 1738175533
transform 1 0 24840 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _0960_
timestamp 1738175533
transform 1 0 25208 0 -1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__nand3_4  _0971_
timestamp 1738175533
transform 1 0 23184 0 1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__dfxtp_2  _1637_
timestamp 1738175533
transform 1 0 25392 0 1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_1  _1672_
timestamp 1738175533
transform 1 0 26864 0 -1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1738175533
transform 1 0 27324 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_281
timestamp 1738175533
transform 1 0 26956 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_286
timestamp 1738175533
transform 1 0 27416 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_276
timestamp 1738175533
transform 1 0 26496 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _0808_
timestamp 1738175533
transform 1 0 28060 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_4  _1069_
timestamp 1738175533
transform -1 0 30912 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _1456_
timestamp 1738175533
transform 1 0 29072 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_292
timestamp 1738175533
transform 1 0 27968 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_302
timestamp 1738175533
transform 1 0 28888 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_300
timestamp 1738175533
transform 1 0 28704 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_307
timestamp 1738175533
transform 1 0 29348 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _0827_
timestamp 1738175533
transform 1 0 31280 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _1574_
timestamp 1738175533
transform 1 0 30636 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1738175533
transform 1 0 29992 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_324
timestamp 1738175533
transform 1 0 30912 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_313
timestamp 1738175533
transform 1 0 29900 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_315
timestamp 1738175533
transform 1 0 30084 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_330
timestamp 1738175533
transform 1 0 31464 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _1760_
timestamp 1738175533
transform 1 0 31832 0 -1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1738175533
transform 1 0 32568 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_335
timestamp 1738175533
transform 1 0 31924 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_341
timestamp 1738175533
transform 1 0 32476 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_343
timestamp 1738175533
transform 1 0 32660 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_355
timestamp 1738175533
transform 1 0 33764 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_354
timestamp 1738175533
transform 1 0 33672 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1738175533
transform -1 0 34316 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1738175533
transform -1 0 34316 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1777_
timestamp 1738175533
transform -1 0 2852 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1738175533
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_19
timestamp 1738175533
transform 1 0 2852 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_23
timestamp 1738175533
transform 1 0 3220 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _0865_
timestamp 1738175533
transform 1 0 5152 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1776_
timestamp 1738175533
transform -1 0 4784 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_40
timestamp 1738175533
transform 1 0 4784 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_47
timestamp 1738175533
transform 1 0 5428 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1269_
timestamp 1738175533
transform 1 0 6808 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1738175533
transform 1 0 6348 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_55
timestamp 1738175533
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_58
timestamp 1738175533
transform 1 0 6440 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_71
timestamp 1738175533
transform 1 0 7636 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__inv_4  _1393_
timestamp 1738175533
transform -1 0 8464 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1590_
timestamp 1738175533
transform 1 0 8832 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_41_80
timestamp 1738175533
transform 1 0 8464 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_93
timestamp 1738175533
transform 1 0 9660 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1738175533
transform -1 0 10304 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1267_
timestamp 1738175533
transform -1 0 12420 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1522_
timestamp 1738175533
transform -1 0 10948 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1738175533
transform 1 0 11592 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_100
timestamp 1738175533
transform 1 0 10304 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_107
timestamp 1738175533
transform 1 0 10948 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_113
timestamp 1738175533
transform 1 0 11500 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_115
timestamp 1738175533
transform 1 0 11684 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_clk_48
timestamp 1738175533
transform -1 0 13892 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1738175533
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_135
timestamp 1738175533
transform 1 0 13524 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_139
timestamp 1738175533
transform 1 0 13892 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1004_
timestamp 1738175533
transform 1 0 16008 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _1073_
timestamp 1738175533
transform -1 0 15640 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_41_147
timestamp 1738175533
transform 1 0 14628 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_158
timestamp 1738175533
transform 1 0 15640 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_166
timestamp 1738175533
transform 1 0 16376 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1005_
timestamp 1738175533
transform 1 0 17296 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1738175533
transform 1 0 16836 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_170
timestamp 1738175533
transform 1 0 16744 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_172
timestamp 1738175533
transform 1 0 16928 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_184
timestamp 1738175533
transform 1 0 18032 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _1729_
timestamp 1738175533
transform 1 0 18860 0 1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_41_192
timestamp 1738175533
transform 1 0 18768 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_213
timestamp 1738175533
transform 1 0 20700 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1738175533
transform 1 0 22632 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1416_
timestamp 1738175533
transform 1 0 21252 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1738175533
transform 1 0 22080 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_223
timestamp 1738175533
transform 1 0 21620 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_227
timestamp 1738175533
transform 1 0 21988 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_229
timestamp 1738175533
transform 1 0 22172 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_233
timestamp 1738175533
transform 1 0 22540 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_237
timestamp 1738175533
transform 1 0 22908 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _0970_
timestamp 1738175533
transform 1 0 23368 0 1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_clk_48
timestamp 1738175533
transform -1 0 25300 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_241
timestamp 1738175533
transform 1 0 23276 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_256
timestamp 1738175533
transform 1 0 24656 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1738175533
transform 1 0 27324 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_263
timestamp 1738175533
transform 1 0 25300 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_275
timestamp 1738175533
transform 1 0 26404 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_283
timestamp 1738175533
transform 1 0 27140 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_286
timestamp 1738175533
transform 1 0 27416 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1457_
timestamp 1738175533
transform 1 0 27968 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_296
timestamp 1738175533
transform 1 0 28336 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_308
timestamp 1738175533
transform 1 0 29440 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0995_
timestamp 1738175533
transform 1 0 29716 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1605_
timestamp 1738175533
transform -1 0 32200 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_318
timestamp 1738175533
transform 1 0 30360 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _0825_
timestamp 1738175533
transform 1 0 33028 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1738175533
transform 1 0 32568 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_338
timestamp 1738175533
transform 1 0 32200 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_343
timestamp 1738175533
transform 1 0 32660 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_352
timestamp 1738175533
transform 1 0 33488 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1738175533
transform -1 0 34316 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0863_
timestamp 1738175533
transform -1 0 2024 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0864_
timestamp 1738175533
transform -1 0 3036 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1738175533
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1738175533
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_10
timestamp 1738175533
transform 1 0 2024 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_21
timestamp 1738175533
transform 1 0 3036 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0866_
timestamp 1738175533
transform 1 0 4508 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1738175533
transform 1 0 3772 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_30
timestamp 1738175533
transform 1 0 3864 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_36
timestamp 1738175533
transform 1 0 4416 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_45
timestamp 1738175533
transform 1 0 5244 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _1676_
timestamp 1738175533
transform -1 0 7452 0 -1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_42_69
timestamp 1738175533
transform 1 0 7452 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1256_
timestamp 1738175533
transform 1 0 7912 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1523_
timestamp 1738175533
transform -1 0 9936 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1738175533
transform 1 0 9016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_73
timestamp 1738175533
transform 1 0 7820 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_78
timestamp 1738175533
transform 1 0 8280 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_87
timestamp 1738175533
transform 1 0 9108 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_2  _1078_
timestamp 1738175533
transform -1 0 11408 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_42_96
timestamp 1738175533
transform 1 0 9936 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_102
timestamp 1738175533
transform 1 0 10488 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_112
timestamp 1738175533
transform 1 0 11408 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1408_
timestamp 1738175533
transform -1 0 13156 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1738175533
transform 1 0 14260 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_120
timestamp 1738175533
transform 1 0 12144 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_131
timestamp 1738175533
transform 1 0 13156 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1767_
timestamp 1738175533
transform 1 0 15180 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_42_144
timestamp 1738175533
transform 1 0 14352 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_152
timestamp 1738175533
transform 1 0 15088 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1766_
timestamp 1738175533
transform -1 0 19044 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_42_169
timestamp 1738175533
transform 1 0 16652 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_177
timestamp 1738175533
transform 1 0 17388 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1738175533
transform 1 0 19504 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_195
timestamp 1738175533
transform 1 0 19044 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_199
timestamp 1738175533
transform 1 0 19412 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_201
timestamp 1738175533
transform 1 0 19596 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_213
timestamp 1738175533
transform 1 0 20700 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_225
timestamp 1738175533
transform 1 0 21804 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_237
timestamp 1738175533
transform 1 0 22908 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_2  _0967_
timestamp 1738175533
transform -1 0 24380 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0969_
timestamp 1738175533
transform -1 0 23552 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1738175533
transform 1 0 24748 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_244
timestamp 1738175533
transform 1 0 23552 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_253
timestamp 1738175533
transform 1 0 24380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_258
timestamp 1738175533
transform 1 0 24840 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1641_
timestamp 1738175533
transform -1 0 26864 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_42_280
timestamp 1738175533
transform 1 0 26864 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _0822_
timestamp 1738175533
transform -1 0 29624 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1455_
timestamp 1738175533
transform 1 0 28152 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_42_292
timestamp 1738175533
transform 1 0 27968 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_299
timestamp 1738175533
transform 1 0 28612 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_4  _0826_
timestamp 1738175533
transform 1 0 30912 0 -1 25568
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1738175533
transform 1 0 29992 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_310
timestamp 1738175533
transform 1 0 29624 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_315
timestamp 1738175533
transform 1 0 30084 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_323
timestamp 1738175533
transform 1 0 30820 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  input9
timestamp 1738175533
transform -1 0 33672 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_42_341
timestamp 1738175533
transform 1 0 32476 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_354
timestamp 1738175533
transform 1 0 33672 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1738175533
transform -1 0 34316 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0849_
timestamp 1738175533
transform 1 0 3036 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1738175533
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1738175533
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_15
timestamp 1738175533
transform 1 0 2484 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0842_
timestamp 1738175533
transform 1 0 4876 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1738175533
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_39
timestamp 1738175533
transform 1 0 4692 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1738175533
transform 1 0 5428 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1580_
timestamp 1738175533
transform -1 0 8004 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1738175533
transform 1 0 6348 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_55
timestamp 1738175533
transform 1 0 6164 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_58
timestamp 1738175533
transform 1 0 6440 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1589_
timestamp 1738175533
transform -1 0 9568 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_43_75
timestamp 1738175533
transform 1 0 8004 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_92
timestamp 1738175533
transform 1 0 9568 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1076_
timestamp 1738175533
transform 1 0 12052 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1449_
timestamp 1738175533
transform -1 0 10580 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1738175533
transform 1 0 11592 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_clk_48
timestamp 1738175533
transform 1 0 10948 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_103
timestamp 1738175533
transform 1 0 10580 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_110
timestamp 1738175533
transform 1 0 11224 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_115
timestamp 1738175533
transform 1 0 11684 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _1656_
timestamp 1738175533
transform 1 0 12788 0 1 25568
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_43_122
timestamp 1738175533
transform 1 0 12328 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_126
timestamp 1738175533
transform 1 0 12696 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1738175533
transform -1 0 16192 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _1397_
timestamp 1738175533
transform -1 0 15548 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_43_148
timestamp 1738175533
transform 1 0 14720 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_157
timestamp 1738175533
transform 1 0 15548 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_164
timestamp 1738175533
transform 1 0 16192 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1001_
timestamp 1738175533
transform 1 0 17296 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1738175533
transform 1 0 16836 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_170
timestamp 1738175533
transform 1 0 16744 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_172
timestamp 1738175533
transform 1 0 16928 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_179
timestamp 1738175533
transform 1 0 17572 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__dfstp_1  _1738_
timestamp 1738175533
transform 1 0 19228 0 1 25568
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_43_191
timestamp 1738175533
transform 1 0 18676 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0981_
timestamp 1738175533
transform 1 0 22816 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1738175533
transform 1 0 22080 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_218
timestamp 1738175533
transform 1 0 21160 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_226
timestamp 1738175533
transform 1 0 21896 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_229
timestamp 1738175533
transform 1 0 22172 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_235
timestamp 1738175533
transform 1 0 22724 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1738175533
transform -1 0 25392 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0955_
timestamp 1738175533
transform 1 0 24288 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_43_242
timestamp 1738175533
transform 1 0 23368 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_250
timestamp 1738175533
transform 1 0 24104 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_257
timestamp 1738175533
transform 1 0 24748 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1299_
timestamp 1738175533
transform 1 0 25852 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1738175533
transform 1 0 27324 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_264
timestamp 1738175533
transform 1 0 25392 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_268
timestamp 1738175533
transform 1 0 25760 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_278
timestamp 1738175533
transform 1 0 26680 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_284
timestamp 1738175533
transform 1 0 27232 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_286
timestamp 1738175533
transform 1 0 27416 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _1671_
timestamp 1738175533
transform 1 0 28152 0 1 25568
box -38 -48 2154 592
use sky130_fd_sc_hd__o21bai_4  _0823_
timestamp 1738175533
transform 1 0 30728 0 1 25568
box -38 -48 1418 592
use sky130_fd_sc_hd__decap_4  FILLER_43_317
timestamp 1738175533
transform 1 0 30268 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_321
timestamp 1738175533
transform 1 0 30636 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _0819_
timestamp 1738175533
transform 1 0 33028 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1738175533
transform 1 0 32568 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_337
timestamp 1738175533
transform 1 0 32108 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_341
timestamp 1738175533
transform 1 0 32476 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_343
timestamp 1738175533
transform 1 0 32660 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_352
timestamp 1738175533
transform 1 0 33488 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1738175533
transform -1 0 34316 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0860_
timestamp 1738175533
transform -1 0 3404 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1738175533
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1738175533
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_15
timestamp 1738175533
transform 1 0 2484 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_19
timestamp 1738175533
transform 1 0 2852 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _0843_
timestamp 1738175533
transform -1 0 5612 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1738175533
transform 1 0 3772 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_25
timestamp 1738175533
transform 1 0 3404 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_30
timestamp 1738175533
transform 1 0 3864 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_38
timestamp 1738175533
transform 1 0 4600 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1579_
timestamp 1738175533
transform -1 0 7912 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_44_49
timestamp 1738175533
transform 1 0 5612 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_61
timestamp 1738175533
transform 1 0 6716 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1294_
timestamp 1738175533
transform 1 0 8280 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1738175533
transform 1 0 9016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_74
timestamp 1738175533
transform 1 0 7912 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_81
timestamp 1738175533
transform 1 0 8556 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_85
timestamp 1738175533
transform 1 0 8924 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_87
timestamp 1738175533
transform 1 0 9108 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_95
timestamp 1738175533
transform 1 0 9844 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_2  _1271_
timestamp 1738175533
transform -1 0 11868 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1563_
timestamp 1738175533
transform 1 0 10028 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_106
timestamp 1738175533
transform 1 0 10856 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_117
timestamp 1738175533
transform 1 0 11868 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1077_
timestamp 1738175533
transform -1 0 13892 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1404_
timestamp 1738175533
transform 1 0 12236 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1738175533
transform 1 0 14260 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_126
timestamp 1738175533
transform 1 0 12696 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_134
timestamp 1738175533
transform 1 0 13432 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_139
timestamp 1738175533
transform 1 0 13892 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_8  _0883_
timestamp 1738175533
transform -1 0 16192 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_44_144
timestamp 1738175533
transform 1 0 14352 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_164
timestamp 1738175533
transform 1 0 16192 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _0818_
timestamp 1738175533
transform -1 0 17296 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_44_168
timestamp 1738175533
transform 1 0 16560 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_176
timestamp 1738175533
transform 1 0 17296 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_188
timestamp 1738175533
transform 1 0 18400 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0987_
timestamp 1738175533
transform 1 0 18676 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__dfstp_1  _1752_
timestamp 1738175533
transform 1 0 20700 0 -1 26656
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1738175533
transform 1 0 19504 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_196
timestamp 1738175533
transform 1 0 19136 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_201
timestamp 1738175533
transform 1 0 19596 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _0983_
timestamp 1738175533
transform -1 0 23460 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_44_234
timestamp 1738175533
transform 1 0 22632 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0959_
timestamp 1738175533
transform -1 0 25668 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0982_
timestamp 1738175533
transform -1 0 24380 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1738175533
transform 1 0 24748 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_243
timestamp 1738175533
transform 1 0 23460 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_247
timestamp 1738175533
transform 1 0 23828 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_253
timestamp 1738175533
transform 1 0 24380 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_258
timestamp 1738175533
transform 1 0 24840 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _1673_
timestamp 1738175533
transform 1 0 26036 0 -1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_44_267
timestamp 1738175533
transform 1 0 25668 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0821_
timestamp 1738175533
transform -1 0 29624 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_44_291
timestamp 1738175533
transform 1 0 27876 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_303
timestamp 1738175533
transform 1 0 28980 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_2  _0824_
timestamp 1738175533
transform 1 0 30728 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1603_
timestamp 1738175533
transform 1 0 31740 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1738175533
transform 1 0 29992 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_310
timestamp 1738175533
transform 1 0 29624 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_315
timestamp 1738175533
transform 1 0 30084 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_321
timestamp 1738175533
transform 1 0 30636 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_329
timestamp 1738175533
transform 1 0 31372 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_349
timestamp 1738175533
transform 1 0 33212 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_357
timestamp 1738175533
transform 1 0 33948 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1738175533
transform -1 0 34316 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1778_
timestamp 1738175533
transform 1 0 1472 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1738175533
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_3
timestamp 1738175533
transform 1 0 1380 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_20
timestamp 1738175533
transform 1 0 2944 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1557_
timestamp 1738175533
transform 1 0 3312 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1785_
timestamp 1738175533
transform 1 0 4508 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_45_33
timestamp 1738175533
transform 1 0 4140 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1575_
timestamp 1738175533
transform 1 0 7452 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1738175533
transform 1 0 6348 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_53
timestamp 1738175533
transform 1 0 5980 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_58
timestamp 1738175533
transform 1 0 6440 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_66
timestamp 1738175533
transform 1 0 7176 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_2  _1295_
timestamp 1738175533
transform 1 0 8648 0 1 26656
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_45_78
timestamp 1738175533
transform 1 0 8280 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_92
timestamp 1738175533
transform 1 0 9568 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1471_
timestamp 1738175533
transform 1 0 10396 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1738175533
transform 1 0 11592 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_100
timestamp 1738175533
transform 1 0 10304 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_107
timestamp 1738175533
transform 1 0 10948 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_113
timestamp 1738175533
transform 1 0 11500 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_115
timestamp 1738175533
transform 1 0 11684 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1075_
timestamp 1738175533
transform -1 0 12512 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1270_
timestamp 1738175533
transform 1 0 13984 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1473_
timestamp 1738175533
transform 1 0 13248 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_clk_48
timestamp 1738175533
transform -1 0 13156 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_124
timestamp 1738175533
transform 1 0 12512 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_131
timestamp 1738175533
transform 1 0 13156 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_136
timestamp 1738175533
transform 1 0 13616 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_143
timestamp 1738175533
transform 1 0 14260 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1608_
timestamp 1738175533
transform 1 0 14996 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_clk_48
timestamp 1738175533
transform 1 0 14628 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_150
timestamp 1738175533
transform 1 0 14904 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _0958_
timestamp 1738175533
transform 1 0 17296 0 1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1738175533
transform 1 0 16836 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_167
timestamp 1738175533
transform 1 0 16468 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_172
timestamp 1738175533
transform 1 0 16928 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_189
timestamp 1738175533
transform 1 0 18492 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1060_
timestamp 1738175533
transform 1 0 20424 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  repeater44
timestamp 1738175533
transform 1 0 18952 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_193
timestamp 1738175533
transform 1 0 18860 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_206
timestamp 1738175533
transform 1 0 20056 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _1041_
timestamp 1738175533
transform 1 0 22540 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1738175533
transform 1 0 22080 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_219
timestamp 1738175533
transform 1 0 21252 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_227
timestamp 1738175533
transform 1 0 21988 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_229
timestamp 1738175533
transform 1 0 22172 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_238
timestamp 1738175533
transform 1 0 23000 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1025_
timestamp 1738175533
transform -1 0 24840 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1040_
timestamp 1738175533
transform -1 0 23644 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_clk_48
timestamp 1738175533
transform -1 0 24288 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_245
timestamp 1738175533
transform 1 0 23644 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_258
timestamp 1738175533
transform 1 0 24840 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1738175533
transform 1 0 27324 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_270
timestamp 1738175533
transform 1 0 25944 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_282
timestamp 1738175533
transform 1 0 27048 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_286
timestamp 1738175533
transform 1 0 27416 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1454_
timestamp 1738175533
transform 1 0 27784 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__buf_8  repeater49
timestamp 1738175533
transform -1 0 30360 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_297
timestamp 1738175533
transform 1 0 28428 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_305
timestamp 1738175533
transform 1 0 29164 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1604_
timestamp 1738175533
transform 1 0 30728 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_45_318
timestamp 1738175533
transform 1 0 30360 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0820_
timestamp 1738175533
transform -1 0 33488 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1738175533
transform 1 0 32568 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_338
timestamp 1738175533
transform 1 0 32200 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_343
timestamp 1738175533
transform 1 0 32660 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_352
timestamp 1738175533
transform 1 0 33488 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1738175533
transform -1 0 34316 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0861_
timestamp 1738175533
transform 1 0 2668 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1738175533
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1738175533
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1738175533
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_15
timestamp 1738175533
transform 1 0 2484 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1738175533
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_15
timestamp 1738175533
transform 1 0 2484 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_23
timestamp 1738175533
transform 1 0 3220 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0845_
timestamp 1738175533
transform 1 0 3496 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1738175533
transform 1 0 3772 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1738175533
transform 1 0 3312 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_28
timestamp 1738175533
transform 1 0 3680 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_30
timestamp 1738175533
transform 1 0 3864 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_30
timestamp 1738175533
transform 1 0 3864 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0833_
timestamp 1738175533
transform 1 0 4232 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1558_
timestamp 1738175533
transform 1 0 4232 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_46_43
timestamp 1738175533
transform 1 0 5060 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_38
timestamp 1738175533
transform 1 0 4600 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0847_
timestamp 1738175533
transform 1 0 5152 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _1643_
timestamp 1738175533
transform -1 0 7544 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1738175533
transform 1 0 6348 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_51
timestamp 1738175533
transform 1 0 5796 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_70
timestamp 1738175533
transform 1 0 7544 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_49
timestamp 1738175533
transform 1 0 5612 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_58
timestamp 1738175533
transform 1 0 6440 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_70
timestamp 1738175533
transform 1 0 7544 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1296_
timestamp 1738175533
transform 1 0 8188 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1461_
timestamp 1738175533
transform 1 0 8096 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_76
timestamp 1738175533
transform 1 0 8096 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_81
timestamp 1738175533
transform 1 0 8556 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1275_
timestamp 1738175533
transform -1 0 10304 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1738175533
transform 1 0 9016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_85
timestamp 1738175533
transform 1 0 8924 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_87
timestamp 1738175533
transform 1 0 9108 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_95
timestamp 1738175533
transform 1 0 9844 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_91
timestamp 1738175533
transform 1 0 9476 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_79
timestamp 1738175533
transform 1 0 8372 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _1272_
timestamp 1738175533
transform 1 0 10028 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1278_
timestamp 1738175533
transform -1 0 11224 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_102
timestamp 1738175533
transform 1 0 10488 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_100
timestamp 1738175533
transform 1 0 10304 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_106
timestamp 1738175533
transform 1 0 10856 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1463_
timestamp 1738175533
transform 1 0 11960 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1465_
timestamp 1738175533
transform 1 0 11316 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1738175533
transform 1 0 11592 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_110
timestamp 1738175533
transform 1 0 11224 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_114
timestamp 1738175533
transform 1 0 11592 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_110
timestamp 1738175533
transform 1 0 11224 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_115
timestamp 1738175533
transform 1 0 11684 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1464_
timestamp 1738175533
transform -1 0 13064 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1549_
timestamp 1738175533
transform 1 0 14168 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1550_
timestamp 1738175533
transform 1 0 13064 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1738175533
transform 1 0 14260 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_121
timestamp 1738175533
transform 1 0 12236 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_129
timestamp 1738175533
transform 1 0 12972 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_139
timestamp 1738175533
transform 1 0 13892 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_130
timestamp 1738175533
transform 1 0 13064 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1548_
timestamp 1738175533
transform 1 0 14720 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_46_144
timestamp 1738175533
transform 1 0 14352 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_157
timestamp 1738175533
transform 1 0 15548 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_151
timestamp 1738175533
transform 1 0 14996 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_163
timestamp 1738175533
transform 1 0 16100 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1061_
timestamp 1738175533
transform 1 0 18492 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1582_
timestamp 1738175533
transform 1 0 17296 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _1737_
timestamp 1738175533
transform 1 0 17204 0 -1 27744
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1738175533
transform 1 0 16836 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_169
timestamp 1738175533
transform 1 0 16652 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_172
timestamp 1738175533
transform 1 0 16928 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_185
timestamp 1738175533
transform 1 0 18124 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_196
timestamp 1738175533
transform 1 0 19136 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_198
timestamp 1738175533
transform 1 0 19320 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1056_
timestamp 1738175533
transform -1 0 20424 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1738175533
transform 1 0 19504 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk_48
timestamp 1738175533
transform -1 0 20240 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_201
timestamp 1738175533
transform 1 0 19596 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_208
timestamp 1738175533
transform 1 0 20240 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_206
timestamp 1738175533
transform 1 0 20056 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _0984_
timestamp 1738175533
transform 1 0 20792 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1057_
timestamp 1738175533
transform 1 0 20700 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_212
timestamp 1738175533
transform 1 0 20608 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_210
timestamp 1738175533
transform 1 0 20424 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1738175533
transform 1 0 21436 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1039_
timestamp 1738175533
transform 1 0 21620 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_217
timestamp 1738175533
transform 1 0 21068 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_217
timestamp 1738175533
transform 1 0 21068 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_224
timestamp 1738175533
transform 1 0 21712 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1034_
timestamp 1738175533
transform 1 0 22908 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1038_
timestamp 1738175533
transform -1 0 22908 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1738175533
transform 1 0 22080 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_227
timestamp 1738175533
transform 1 0 21988 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_229
timestamp 1738175533
transform 1 0 22172 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_237
timestamp 1738175533
transform 1 0 22908 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_241
timestamp 1738175533
transform 1 0 23276 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_245
timestamp 1738175533
transform 1 0 23644 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_1  _1093_
timestamp 1738175533
transform 1 0 23736 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_249
timestamp 1738175533
transform 1 0 24012 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_252
timestamp 1738175533
transform 1 0 24288 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1027_
timestamp 1738175533
transform -1 0 25024 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1738175533
transform 1 0 24748 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_clk_48
timestamp 1738175533
transform -1 0 24656 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_256
timestamp 1738175533
transform 1 0 24656 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_258
timestamp 1738175533
transform 1 0 24840 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1026_
timestamp 1738175533
transform -1 0 25484 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_260
timestamp 1738175533
transform 1 0 25024 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1030_
timestamp 1738175533
transform 1 0 26312 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1031_
timestamp 1738175533
transform 1 0 25392 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1738175533
transform 1 0 27324 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1738175533
transform 1 0 25484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1738175533
transform 1 0 26588 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_270
timestamp 1738175533
transform 1 0 25944 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_277
timestamp 1738175533
transform 1 0 26588 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_286
timestamp 1738175533
transform 1 0 27416 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0830_
timestamp 1738175533
transform 1 0 28796 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _1786_
timestamp 1738175533
transform 1 0 28428 0 1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1738175533
transform 1 0 27692 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_308
timestamp 1738175533
transform 1 0 29440 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_47_294
timestamp 1738175533
transform 1 0 28152 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0810_
timestamp 1738175533
transform 1 0 31464 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0829_
timestamp 1738175533
transform -1 0 31096 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _1602_
timestamp 1738175533
transform -1 0 32016 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1738175533
transform 1 0 29992 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_315
timestamp 1738175533
transform 1 0 30084 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_319
timestamp 1738175533
transform 1 0 30452 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_317
timestamp 1738175533
transform 1 0 30268 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_326
timestamp 1738175533
transform 1 0 31096 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1409_
timestamp 1738175533
transform -1 0 32844 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1738175533
transform 1 0 32568 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_336
timestamp 1738175533
transform 1 0 32016 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1738175533
transform 1 0 32844 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_357
timestamp 1738175533
transform 1 0 33948 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_334
timestamp 1738175533
transform 1 0 31832 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_343
timestamp 1738175533
transform 1 0 32660 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_355
timestamp 1738175533
transform 1 0 33764 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1738175533
transform -1 0 34316 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1738175533
transform -1 0 34316 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1779_
timestamp 1738175533
transform 1 0 1748 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1738175533
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1738175533
transform 1 0 1380 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_23
timestamp 1738175533
transform 1 0 3220 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1784_
timestamp 1738175533
transform 1 0 4784 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1738175533
transform 1 0 3772 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_30
timestamp 1738175533
transform 1 0 3864 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_38
timestamp 1738175533
transform 1 0 4600 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1556_
timestamp 1738175533
transform 1 0 6624 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_48_56
timestamp 1738175533
transform 1 0 6256 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_69
timestamp 1738175533
transform 1 0 7452 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1470_
timestamp 1738175533
transform 1 0 8372 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1547_
timestamp 1738175533
transform -1 0 10304 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1738175533
transform 1 0 9016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_77
timestamp 1738175533
transform 1 0 8188 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_82
timestamp 1738175533
transform 1 0 8648 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_87
timestamp 1738175533
transform 1 0 9108 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1649_
timestamp 1738175533
transform 1 0 10948 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_48_100
timestamp 1738175533
transform 1 0 10304 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_106
timestamp 1738175533
transform 1 0 10856 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1277_
timestamp 1738175533
transform -1 0 13064 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1472_
timestamp 1738175533
transform 1 0 13616 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1738175533
transform 1 0 14260 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_123
timestamp 1738175533
transform 1 0 12420 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_130
timestamp 1738175533
transform 1 0 13064 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_139
timestamp 1738175533
transform 1 0 13892 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1594_
timestamp 1738175533
transform 1 0 14720 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_48_144
timestamp 1738175533
transform 1 0 14352 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_157
timestamp 1738175533
transform 1 0 15548 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_165
timestamp 1738175533
transform 1 0 16284 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1388_
timestamp 1738175533
transform 1 0 16560 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_48_173
timestamp 1738175533
transform 1 0 17020 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_185
timestamp 1738175533
transform 1 0 18124 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _0989_
timestamp 1738175533
transform -1 0 19136 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _0993_
timestamp 1738175533
transform 1 0 19964 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1738175533
transform 1 0 19504 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_191
timestamp 1738175533
transform 1 0 18676 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_196
timestamp 1738175533
transform 1 0 19136 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_201
timestamp 1738175533
transform 1 0 19596 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_209
timestamp 1738175533
transform 1 0 20332 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1058_
timestamp 1738175533
transform -1 0 22264 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _1059_
timestamp 1738175533
transform 1 0 20884 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_48_220
timestamp 1738175533
transform 1 0 21344 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_226
timestamp 1738175533
transform 1 0 21896 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_230
timestamp 1738175533
transform 1 0 22264 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_1  _1028_
timestamp 1738175533
transform 1 0 25208 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1037_
timestamp 1738175533
transform 1 0 23644 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1738175533
transform 1 0 24748 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_242
timestamp 1738175533
transform 1 0 23368 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_252
timestamp 1738175533
transform 1 0 24288 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_256
timestamp 1738175533
transform 1 0 24656 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_258
timestamp 1738175533
transform 1 0 24840 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _1755_
timestamp 1738175533
transform -1 0 27968 0 -1 28832
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_48_267
timestamp 1738175533
transform 1 0 25668 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0816_
timestamp 1738175533
transform 1 0 28796 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_48_292
timestamp 1738175533
transform 1 0 27968 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_300
timestamp 1738175533
transform 1 0 28704 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__or3b_4  _1412_
timestamp 1738175533
transform 1 0 30452 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1738175533
transform 1 0 29992 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_310
timestamp 1738175533
transform 1 0 29624 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_315
timestamp 1738175533
transform 1 0 30084 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_328
timestamp 1738175533
transform 1 0 31280 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1601_
timestamp 1738175533
transform 1 0 32108 0 -1 28832
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_48_336
timestamp 1738175533
transform 1 0 32016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_354
timestamp 1738175533
transform 1 0 33672 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1738175533
transform -1 0 34316 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0859_
timestamp 1738175533
transform 1 0 3036 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1738175533
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1738175533
transform -1 0 2024 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 1738175533
transform 1 0 1380 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_10
timestamp 1738175533
transform 1 0 2024 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_18
timestamp 1738175533
transform 1 0 2760 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0848_
timestamp 1738175533
transform 1 0 5060 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0858_
timestamp 1738175533
transform -1 0 4508 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_49_28
timestamp 1738175533
transform 1 0 3680 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_37
timestamp 1738175533
transform 1 0 4508 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1545_
timestamp 1738175533
transform -1 0 8096 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1738175533
transform 1 0 6348 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_50
timestamp 1738175533
transform 1 0 5704 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_56
timestamp 1738175533
transform 1 0 6256 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_58
timestamp 1738175533
transform 1 0 6440 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_66
timestamp 1738175533
transform 1 0 7176 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1276_
timestamp 1738175533
transform 1 0 9660 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1577_
timestamp 1738175533
transform 1 0 8464 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_49_76
timestamp 1738175533
transform 1 0 8096 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_89
timestamp 1738175533
transform 1 0 9292 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1274_
timestamp 1738175533
transform -1 0 10764 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1738175533
transform 1 0 11592 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_97
timestamp 1738175533
transform 1 0 10028 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_101
timestamp 1738175533
transform 1 0 10396 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_105
timestamp 1738175533
transform 1 0 10764 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_113
timestamp 1738175533
transform 1 0 11500 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_115
timestamp 1738175533
transform 1 0 11684 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1542_
timestamp 1738175533
transform 1 0 12696 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1595_
timestamp 1738175533
transform -1 0 15088 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_clk_48
timestamp 1738175533
transform 1 0 12420 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_135
timestamp 1738175533
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_152
timestamp 1738175533
transform 1 0 15088 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_164
timestamp 1738175533
transform 1 0 16192 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1054_
timestamp 1738175533
transform 1 0 18308 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__nor2b_1  _1389_
timestamp 1738175533
transform 1 0 17296 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1738175533
transform 1 0 16836 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_170
timestamp 1738175533
transform 1 0 16744 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_172
timestamp 1738175533
transform 1 0 16928 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_181
timestamp 1738175533
transform 1 0 17756 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0986_
timestamp 1738175533
transform -1 0 20608 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_196
timestamp 1738175533
transform 1 0 19136 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_208
timestamp 1738175533
transform 1 0 20240 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_212
timestamp 1738175533
transform 1 0 20608 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1738175533
transform 1 0 22080 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_224
timestamp 1738175533
transform 1 0 21712 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_229
timestamp 1738175533
transform 1 0 22172 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1036_
timestamp 1738175533
transform 1 0 24196 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1091_
timestamp 1738175533
transform 1 0 25116 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_clk_48
timestamp 1738175533
transform 1 0 23368 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_241
timestamp 1738175533
transform 1 0 23276 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_245
timestamp 1738175533
transform 1 0 23644 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_254
timestamp 1738175533
transform 1 0 24472 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_260
timestamp 1738175533
transform 1 0 25024 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1738175533
transform 1 0 27324 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_clk_48
timestamp 1738175533
transform -1 0 26588 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_266
timestamp 1738175533
transform 1 0 25576 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_277
timestamp 1738175533
transform 1 0 26588 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_286
timestamp 1738175533
transform 1 0 27416 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _1787_
timestamp 1738175533
transform 1 0 27968 0 1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  _0815_
timestamp 1738175533
transform 1 0 30636 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_49_312
timestamp 1738175533
transform 1 0 29808 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_320
timestamp 1738175533
transform 1 0 30544 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_330
timestamp 1738175533
transform 1 0 31464 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1738175533
transform 1 0 32568 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1738175533
transform 1 0 33396 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_343
timestamp 1738175533
transform 1 0 32660 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_354
timestamp 1738175533
transform 1 0 33672 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1738175533
transform -1 0 34316 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0856_
timestamp 1738175533
transform -1 0 3404 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1738175533
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1738175533
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_15
timestamp 1738175533
transform 1 0 2484 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_19
timestamp 1738175533
transform 1 0 2852 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1551_
timestamp 1738175533
transform 1 0 4232 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1738175533
transform 1 0 3772 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_25
timestamp 1738175533
transform 1 0 3404 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_30
timestamp 1738175533
transform 1 0 3864 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_43
timestamp 1738175533
transform 1 0 5060 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_47
timestamp 1738175533
transform 1 0 5428 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _0835_
timestamp 1738175533
transform -1 0 5980 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1546_
timestamp 1738175533
transform -1 0 8188 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1738175533
transform 1 0 5980 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_65
timestamp 1738175533
transform 1 0 7084 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1281_
timestamp 1738175533
transform 1 0 9476 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1738175533
transform 1 0 9016 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_77
timestamp 1738175533
transform 1 0 8188 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_85
timestamp 1738175533
transform 1 0 8924 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_87
timestamp 1738175533
transform 1 0 9108 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_95
timestamp 1738175533
transform 1 0 9844 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1280_
timestamp 1738175533
transform 1 0 10212 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1544_
timestamp 1738175533
transform 1 0 10948 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_50_102
timestamp 1738175533
transform 1 0 10488 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_106
timestamp 1738175533
transform 1 0 10856 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_116
timestamp 1738175533
transform 1 0 11776 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1543_
timestamp 1738175533
transform 1 0 12144 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1738175533
transform 1 0 14260 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_129
timestamp 1738175533
transform 1 0 12972 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1738175533
transform 1 0 14076 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1607_
timestamp 1738175533
transform -1 0 16744 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_clk_48
timestamp 1738175533
transform -1 0 14996 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_144
timestamp 1738175533
transform 1 0 14352 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_151
timestamp 1738175533
transform 1 0 14996 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _1741_
timestamp 1738175533
transform 1 0 17204 0 -1 29920
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_50_170
timestamp 1738175533
transform 1 0 16744 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_174
timestamp 1738175533
transform 1 0 17112 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1738175533
transform 1 0 19504 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_196
timestamp 1738175533
transform 1 0 19136 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_201
timestamp 1738175533
transform 1 0 19596 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_213
timestamp 1738175533
transform 1 0 20700 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _1739_
timestamp 1738175533
transform 1 0 21068 0 -1 29920
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_50_238
timestamp 1738175533
transform 1 0 23000 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1738175533
transform 1 0 25208 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1738175533
transform 1 0 24748 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_250
timestamp 1738175533
transform 1 0 24104 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_256
timestamp 1738175533
transform 1 0 24656 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_258
timestamp 1738175533
transform 1 0 24840 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _1092_
timestamp 1738175533
transform -1 0 26404 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_265
timestamp 1738175533
transform 1 0 25484 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_275
timestamp 1738175533
transform 1 0 26404 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__nor3_4  _1415_
timestamp 1738175533
transform -1 0 28888 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_50_287
timestamp 1738175533
transform 1 0 27508 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_302
timestamp 1738175533
transform 1 0 28888 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _1788_
timestamp 1738175533
transform 1 0 30636 0 -1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1738175533
transform 1 0 29992 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_315
timestamp 1738175533
transform 1 0 30084 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_341
timestamp 1738175533
transform 1 0 32476 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_353
timestamp 1738175533
transform 1 0 33580 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_357
timestamp 1738175533
transform 1 0 33948 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1738175533
transform -1 0 34316 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1780_
timestamp 1738175533
transform 1 0 1380 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1738175533
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_19
timestamp 1738175533
transform 1 0 2852 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_4  _0834_
timestamp 1738175533
transform 1 0 3680 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_51_27
timestamp 1738175533
transform 1 0 3588 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_41
timestamp 1738175533
transform 1 0 4876 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1555_
timestamp 1738175533
transform 1 0 6808 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1738175533
transform 1 0 6348 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_53
timestamp 1738175533
transform 1 0 5980 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_58
timestamp 1738175533
transform 1 0 6440 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_71
timestamp 1738175533
transform 1 0 7636 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1279_
timestamp 1738175533
transform 1 0 8740 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_86
timestamp 1738175533
transform 1 0 9016 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_94
timestamp 1738175533
transform 1 0 9752 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _1289_
timestamp 1738175533
transform -1 0 10856 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1290_
timestamp 1738175533
transform 1 0 9936 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1738175533
transform 1 0 11592 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_clk_48
timestamp 1738175533
transform 1 0 11224 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_99
timestamp 1738175533
transform 1 0 10212 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_106
timestamp 1738175533
transform 1 0 10856 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_113
timestamp 1738175533
transform 1 0 11500 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_115
timestamp 1738175533
transform 1 0 11684 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1292_
timestamp 1738175533
transform -1 0 13340 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1541_
timestamp 1738175533
transform 1 0 13708 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_51_127
timestamp 1738175533
transform 1 0 12788 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_133
timestamp 1738175533
transform 1 0 13340 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1293_
timestamp 1738175533
transform 1 0 14904 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_146
timestamp 1738175533
transform 1 0 14536 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_154
timestamp 1738175533
transform 1 0 15272 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_166
timestamp 1738175533
transform 1 0 16376 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1053_
timestamp 1738175533
transform 1 0 18216 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1738175533
transform 1 0 16836 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_170
timestamp 1738175533
transform 1 0 16744 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_172
timestamp 1738175533
transform 1 0 16928 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_184
timestamp 1738175533
transform 1 0 18032 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_1  _1740_
timestamp 1738175533
transform -1 0 21528 0 1 29920
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_51_195
timestamp 1738175533
transform 1 0 19044 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__dfstp_1  _1753_
timestamp 1738175533
transform 1 0 22632 0 1 29920
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1738175533
transform 1 0 22080 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_222
timestamp 1738175533
transform 1 0 21528 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_229
timestamp 1738175533
transform 1 0 22172 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_233
timestamp 1738175533
transform 1 0 22540 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_255
timestamp 1738175533
transform 1 0 24564 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1022_
timestamp 1738175533
transform 1 0 26036 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1052_
timestamp 1738175533
transform 1 0 25300 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1738175533
transform 1 0 27324 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_267
timestamp 1738175533
transform 1 0 25668 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_280
timestamp 1738175533
transform 1 0 26864 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_284
timestamp 1738175533
transform 1 0 27232 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_286
timestamp 1738175533
transform 1 0 27416 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3b_4  _1414_
timestamp 1738175533
transform 1 0 29072 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_51_298
timestamp 1738175533
transform 1 0 28520 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_320
timestamp 1738175533
transform 1 0 30544 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_332
timestamp 1738175533
transform 1 0 31648 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1738175533
transform 1 0 32568 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_340
timestamp 1738175533
transform 1 0 32384 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_343
timestamp 1738175533
transform 1 0 32660 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_355
timestamp 1738175533
transform 1 0 33764 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1738175533
transform -1 0 34316 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0857_
timestamp 1738175533
transform 1 0 2760 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1738175533
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1738175533
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1738175533
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_15
timestamp 1738175533
transform 1 0 2484 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1738175533
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1738175533
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3_4  _0837_
timestamp 1738175533
transform -1 0 6256 0 -1 31008
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _1552_
timestamp 1738175533
transform 1 0 3588 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1738175533
transform 1 0 3772 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_25
timestamp 1738175533
transform 1 0 3404 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_30
timestamp 1738175533
transform 1 0 3864 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_36
timestamp 1738175533
transform 1 0 4416 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _0836_
timestamp 1738175533
transform -1 0 5980 0 1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0850_
timestamp 1738175533
transform 1 0 6808 0 1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0851_
timestamp 1738175533
transform 1 0 6624 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1738175533
transform 1 0 6348 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_56
timestamp 1738175533
transform 1 0 6256 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_67
timestamp 1738175533
transform 1 0 7268 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_53
timestamp 1738175533
transform 1 0 5980 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_58
timestamp 1738175533
transform 1 0 6440 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_67
timestamp 1738175533
transform 1 0 7268 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1648_
timestamp 1738175533
transform -1 0 9568 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1738175533
transform 1 0 9016 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_79
timestamp 1738175533
transform 1 0 8372 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_85
timestamp 1738175533
transform 1 0 8924 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_87
timestamp 1738175533
transform 1 0 9108 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_75
timestamp 1738175533
transform 1 0 8004 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_92
timestamp 1738175533
transform 1 0 9568 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1288_
timestamp 1738175533
transform -1 0 10396 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1645_
timestamp 1738175533
transform 1 0 10212 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1738175533
transform 1 0 11592 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_115
timestamp 1738175533
transform 1 0 11684 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_101
timestamp 1738175533
transform 1 0 10396 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_113
timestamp 1738175533
transform 1 0 11500 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_115
timestamp 1738175533
transform 1 0 11684 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1462_
timestamp 1738175533
transform -1 0 13984 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1585_
timestamp 1738175533
transform 1 0 12420 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1586_
timestamp 1738175533
transform -1 0 13156 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1738175533
transform 1 0 14260 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_132
timestamp 1738175533
transform 1 0 13248 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_140
timestamp 1738175533
transform 1 0 13984 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_121
timestamp 1738175533
transform 1 0 12236 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_131
timestamp 1738175533
transform 1 0 13156 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_140
timestamp 1738175533
transform 1 0 13984 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1291_
timestamp 1738175533
transform 1 0 14720 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1644_
timestamp 1738175533
transform -1 0 15824 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _1742_
timestamp 1738175533
transform 1 0 16100 0 -1 31008
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_52_144
timestamp 1738175533
transform 1 0 14352 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_151
timestamp 1738175533
transform 1 0 14996 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_160
timestamp 1738175533
transform 1 0 15824 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1051_
timestamp 1738175533
transform 1 0 17480 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1738175533
transform 1 0 16836 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_184
timestamp 1738175533
transform 1 0 18032 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_168
timestamp 1738175533
transform 1 0 16560 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_172
timestamp 1738175533
transform 1 0 16928 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_187
timestamp 1738175533
transform 1 0 18308 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0988_
timestamp 1738175533
transform 1 0 18676 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1055_
timestamp 1738175533
transform 1 0 20148 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1738175533
transform 1 0 19504 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_196
timestamp 1738175533
transform 1 0 19136 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_201
timestamp 1738175533
transform 1 0 19596 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_200
timestamp 1738175533
transform 1 0 19504 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_212
timestamp 1738175533
transform 1 0 20608 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1020_
timestamp 1738175533
transform 1 0 22816 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1045_
timestamp 1738175533
transform -1 0 22908 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1738175533
transform 1 0 22080 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_216
timestamp 1738175533
transform 1 0 20976 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_228
timestamp 1738175533
transform 1 0 22080 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_224
timestamp 1738175533
transform 1 0 21712 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_229
timestamp 1738175533
transform 1 0 22172 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_237
timestamp 1738175533
transform 1 0 22908 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1032_
timestamp 1738175533
transform 1 0 23552 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _1754_
timestamp 1738175533
transform 1 0 23552 0 1 31008
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1738175533
transform 1 0 24748 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_240
timestamp 1738175533
transform 1 0 23184 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_253
timestamp 1738175533
transform 1 0 24380 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_258
timestamp 1738175533
transform 1 0 24840 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_243
timestamp 1738175533
transform 1 0 23460 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _1756_
timestamp 1738175533
transform -1 0 27784 0 -1 31008
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1738175533
transform 1 0 27324 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_266
timestamp 1738175533
transform 1 0 25576 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_265
timestamp 1738175533
transform 1 0 25484 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_277
timestamp 1738175533
transform 1 0 26588 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_286
timestamp 1738175533
transform 1 0 27416 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _1792_
timestamp 1738175533
transform 1 0 27784 0 1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_52_290
timestamp 1738175533
transform 1 0 27784 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_302
timestamp 1738175533
transform 1 0 28888 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0814_
timestamp 1738175533
transform 1 0 30820 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _1789_
timestamp 1738175533
transform 1 0 30728 0 -1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1738175533
transform 1 0 29992 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_315
timestamp 1738175533
transform 1 0 30084 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_321
timestamp 1738175533
transform 1 0 30636 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_310
timestamp 1738175533
transform 1 0 29624 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_322
timestamp 1738175533
transform 1 0 30728 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_332
timestamp 1738175533
transform 1 0 31648 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1738175533
transform 1 0 32568 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_342
timestamp 1738175533
transform 1 0 32568 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_354
timestamp 1738175533
transform 1 0 33672 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_340
timestamp 1738175533
transform 1 0 32384 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_343
timestamp 1738175533
transform 1 0 32660 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_355
timestamp 1738175533
transform 1 0 33764 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1738175533
transform -1 0 34316 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1738175533
transform -1 0 34316 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0854_
timestamp 1738175533
transform 1 0 2944 0 -1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1738175533
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1738175533
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_15
timestamp 1738175533
transform 1 0 2484 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_19
timestamp 1738175533
transform 1 0 2852 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _0852_
timestamp 1738175533
transform 1 0 4324 0 -1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0853_
timestamp 1738175533
transform -1 0 5796 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1738175533
transform 1 0 3772 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_25
timestamp 1738175533
transform 1 0 3404 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_30
timestamp 1738175533
transform 1 0 3864 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_34
timestamp 1738175533
transform 1 0 4232 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_40
timestamp 1738175533
transform 1 0 4784 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1783_
timestamp 1738175533
transform 1 0 6440 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_54_51
timestamp 1738175533
transform 1 0 5796 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_57
timestamp 1738175533
transform 1 0 6348 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1398_
timestamp 1738175533
transform -1 0 9752 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1738175533
transform 1 0 9016 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_74
timestamp 1738175533
transform 1 0 7912 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_87
timestamp 1738175533
transform 1 0 9108 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_94
timestamp 1738175533
transform 1 0 9752 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1283_
timestamp 1738175533
transform 1 0 10120 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_101
timestamp 1738175533
transform 1 0 10396 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_113
timestamp 1738175533
transform 1 0 11500 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1467_
timestamp 1738175533
transform 1 0 12328 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1468_
timestamp 1738175533
transform -1 0 13248 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1738175533
transform 1 0 14260 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_121
timestamp 1738175533
transform 1 0 12236 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_125
timestamp 1738175533
transform 1 0 12604 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_132
timestamp 1738175533
transform 1 0 13248 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_140
timestamp 1738175533
transform 1 0 13984 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1581_
timestamp 1738175533
transform -1 0 15548 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _1743_
timestamp 1738175533
transform 1 0 16192 0 -1 32096
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_54_144
timestamp 1738175533
transform 1 0 14352 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_157
timestamp 1738175533
transform 1 0 15548 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_163
timestamp 1738175533
transform 1 0 16100 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_185
timestamp 1738175533
transform 1 0 18124 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1047_
timestamp 1738175533
transform 1 0 19964 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1738175533
transform 1 0 19504 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_197
timestamp 1738175533
transform 1 0 19228 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_201
timestamp 1738175533
transform 1 0 19596 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_214
timestamp 1738175533
transform 1 0 20792 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__dfstp_1  _1751_
timestamp 1738175533
transform -1 0 23552 0 -1 32096
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_54_222
timestamp 1738175533
transform 1 0 21528 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1738175533
transform 1 0 24748 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_244
timestamp 1738175533
transform 1 0 23552 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_256
timestamp 1738175533
transform 1 0 24656 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_258
timestamp 1738175533
transform 1 0 24840 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__dfstp_1  _1757_
timestamp 1738175533
transform 1 0 25484 0 -1 32096
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_54_264
timestamp 1738175533
transform 1 0 25392 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_286
timestamp 1738175533
transform 1 0 27416 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0811_
timestamp 1738175533
transform 1 0 28612 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_54_298
timestamp 1738175533
transform 1 0 28520 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_308
timestamp 1738175533
transform 1 0 29440 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0813_
timestamp 1738175533
transform 1 0 30452 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1413_
timestamp 1738175533
transform -1 0 32200 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1738175533
transform 1 0 29992 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_315
timestamp 1738175533
transform 1 0 30084 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_328
timestamp 1738175533
transform 1 0 31280 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_338
timestamp 1738175533
transform 1 0 32200 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_350
timestamp 1738175533
transform 1 0 33304 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1738175533
transform -1 0 34316 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1781_
timestamp 1738175533
transform -1 0 3956 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1738175533
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1738175533
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1553_
timestamp 1738175533
transform 1 0 5060 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_55_31
timestamp 1738175533
transform 1 0 3956 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1554_
timestamp 1738175533
transform 1 0 6900 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1738175533
transform 1 0 6348 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1738175533
transform 1 0 5888 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_56
timestamp 1738175533
transform 1 0 6256 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_58
timestamp 1738175533
transform 1 0 6440 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_62
timestamp 1738175533
transform 1 0 6808 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_1  _1287_
timestamp 1738175533
transform 1 0 8280 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1466_
timestamp 1738175533
transform 1 0 9016 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1647_
timestamp 1738175533
transform 1 0 9752 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_55_72
timestamp 1738175533
transform 1 0 7728 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_82
timestamp 1738175533
transform 1 0 8648 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_89
timestamp 1738175533
transform 1 0 9292 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_93
timestamp 1738175533
transform 1 0 9660 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1738175533
transform 1 0 11592 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_110
timestamp 1738175533
transform 1 0 11224 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_115
timestamp 1738175533
transform 1 0 11684 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1576_
timestamp 1738175533
transform -1 0 13156 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1587_
timestamp 1738175533
transform 1 0 13524 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_55_121
timestamp 1738175533
transform 1 0 12236 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_131
timestamp 1738175533
transform 1 0 13156 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1539_
timestamp 1738175533
transform 1 0 14812 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_55_144
timestamp 1738175533
transform 1 0 14352 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_148
timestamp 1738175533
transform 1 0 14720 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_158
timestamp 1738175533
transform 1 0 15640 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1050_
timestamp 1738175533
transform 1 0 17940 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1738175533
transform 1 0 16836 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_170
timestamp 1738175533
transform 1 0 16744 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_172
timestamp 1738175533
transform 1 0 16928 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_180
timestamp 1738175533
transform 1 0 17664 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0992_
timestamp 1738175533
transform -1 0 19412 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _1747_
timestamp 1738175533
transform 1 0 19780 0 1 32096
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_55_192
timestamp 1738175533
transform 1 0 18768 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_199
timestamp 1738175533
transform 1 0 19412 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1042_
timestamp 1738175533
transform -1 0 23368 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1738175533
transform 1 0 22080 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_224
timestamp 1738175533
transform 1 0 21712 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_229
timestamp 1738175533
transform 1 0 22172 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1043_
timestamp 1738175533
transform -1 0 24840 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_55_242
timestamp 1738175533
transform 1 0 23368 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_248
timestamp 1738175533
transform 1 0 23920 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_258
timestamp 1738175533
transform 1 0 24840 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1021_
timestamp 1738175533
transform 1 0 25852 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1738175533
transform 1 0 27324 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_266
timestamp 1738175533
transform 1 0 25576 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_278
timestamp 1738175533
transform 1 0 26680 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_284
timestamp 1738175533
transform 1 0 27232 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_286
timestamp 1738175533
transform 1 0 27416 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0812_
timestamp 1738175533
transform 1 0 28888 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_55_298
timestamp 1738175533
transform 1 0 28520 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _1790_
timestamp 1738175533
transform 1 0 30084 0 1 32096
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_55_311
timestamp 1738175533
transform 1 0 29716 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1738175533
transform 1 0 32568 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_335
timestamp 1738175533
transform 1 0 31924 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_341
timestamp 1738175533
transform 1 0 32476 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_343
timestamp 1738175533
transform 1 0 32660 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_355
timestamp 1738175533
transform 1 0 33764 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1738175533
transform -1 0 34316 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1738175533
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1738175533
transform 1 0 1380 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_6
timestamp 1738175533
transform 1 0 1656 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_18
timestamp 1738175533
transform 1 0 2760 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1782_
timestamp 1738175533
transform -1 0 5980 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1738175533
transform 1 0 3772 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_26
timestamp 1738175533
transform 1 0 3496 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_30
timestamp 1738175533
transform 1 0 3864 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_36
timestamp 1738175533
transform 1 0 4416 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1646_
timestamp 1738175533
transform -1 0 8004 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_56_53
timestamp 1738175533
transform 1 0 5980 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1284_
timestamp 1738175533
transform 1 0 9568 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1285_
timestamp 1738175533
transform 1 0 8372 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1738175533
transform 1 0 9016 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_75
timestamp 1738175533
transform 1 0 8004 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_82
timestamp 1738175533
transform 1 0 8648 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_87
timestamp 1738175533
transform 1 0 9108 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_91
timestamp 1738175533
transform 1 0 9476 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1297_
timestamp 1738175533
transform -1 0 10764 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_98
timestamp 1738175533
transform 1 0 10120 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_105
timestamp 1738175533
transform 1 0 10764 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_117
timestamp 1738175533
transform 1 0 11868 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1588_
timestamp 1738175533
transform 1 0 12420 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1738175533
transform 1 0 14260 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_132
timestamp 1738175533
transform 1 0 13248 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_140
timestamp 1738175533
transform 1 0 13984 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1540_
timestamp 1738175533
transform 1 0 14720 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _1744_
timestamp 1738175533
transform 1 0 16376 0 -1 33184
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_56_144
timestamp 1738175533
transform 1 0 14352 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_157
timestamp 1738175533
transform 1 0 15548 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_165
timestamp 1738175533
transform 1 0 16284 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_187
timestamp 1738175533
transform 1 0 18308 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _0991_
timestamp 1738175533
transform 1 0 19964 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1738175533
transform 1 0 19504 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_199
timestamp 1738175533
transform 1 0 19412 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_201
timestamp 1738175533
transform 1 0 19596 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_214
timestamp 1738175533
transform 1 0 20792 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _0990_
timestamp 1738175533
transform -1 0 23644 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_56_226
timestamp 1738175533
transform 1 0 21896 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_234
timestamp 1738175533
transform 1 0 22632 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1738175533
transform 1 0 24748 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_245
timestamp 1738175533
transform 1 0 23644 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_258
timestamp 1738175533
transform 1 0 24840 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_270
timestamp 1738175533
transform 1 0 25944 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_282
timestamp 1738175533
transform 1 0 27048 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_294
timestamp 1738175533
transform 1 0 28152 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_306
timestamp 1738175533
transform 1 0 29256 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1738175533
transform 1 0 29992 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_315
timestamp 1738175533
transform 1 0 30084 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_327
timestamp 1738175533
transform 1 0 31188 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1469_
timestamp 1738175533
transform 1 0 33396 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_339
timestamp 1738175533
transform 1 0 32292 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_354
timestamp 1738175533
transform 1 0 33672 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1738175533
transform -1 0 34316 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1738175533
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1738175533
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_15
timestamp 1738175533
transform 1 0 2484 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_23
timestamp 1738175533
transform 1 0 3220 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0855_
timestamp 1738175533
transform 1 0 3496 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_57_33
timestamp 1738175533
transform 1 0 4140 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_45
timestamp 1738175533
transform 1 0 5244 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1597_
timestamp 1738175533
transform -1 0 8280 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1738175533
transform 1 0 6348 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_58
timestamp 1738175533
transform 1 0 6440 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_66
timestamp 1738175533
transform 1 0 7176 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_2  _1286_
timestamp 1738175533
transform 1 0 8648 0 1 33184
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_57_78
timestamp 1738175533
transform 1 0 8280 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_92
timestamp 1738175533
transform 1 0 9568 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1273_
timestamp 1738175533
transform -1 0 10672 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1592_
timestamp 1738175533
transform -1 0 12880 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1738175533
transform 1 0 11592 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_104
timestamp 1738175533
transform 1 0 10672 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_112
timestamp 1738175533
transform 1 0 11408 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_115
timestamp 1738175533
transform 1 0 11684 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1459_
timestamp 1738175533
transform 1 0 13248 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_128
timestamp 1738175533
transform 1 0 12880 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_135
timestamp 1738175533
transform 1 0 13524 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_143
timestamp 1738175533
transform 1 0 14260 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _1659_
timestamp 1738175533
transform 1 0 14352 0 1 33184
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_57_164
timestamp 1738175533
transform 1 0 16192 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1049_
timestamp 1738175533
transform 1 0 18124 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1738175533
transform 1 0 16836 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_170
timestamp 1738175533
transform 1 0 16744 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_172
timestamp 1738175533
transform 1 0 16928 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_184
timestamp 1738175533
transform 1 0 18032 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1048_
timestamp 1738175533
transform 1 0 19412 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_57_194
timestamp 1738175533
transform 1 0 18952 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_198
timestamp 1738175533
transform 1 0 19320 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_208
timestamp 1738175533
transform 1 0 20240 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_214
timestamp 1738175533
transform 1 0 20792 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1046_
timestamp 1738175533
transform -1 0 21712 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1738175533
transform 1 0 22080 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_224
timestamp 1738175533
transform 1 0 21712 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_229
timestamp 1738175533
transform 1 0 22172 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__dfstp_1  _1750_
timestamp 1738175533
transform -1 0 25760 0 1 33184
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_57_241
timestamp 1738175533
transform 1 0 23276 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1738175533
transform 1 0 27324 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_268
timestamp 1738175533
transform 1 0 25760 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_280
timestamp 1738175533
transform 1 0 26864 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_284
timestamp 1738175533
transform 1 0 27232 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_286
timestamp 1738175533
transform 1 0 27416 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _1791_
timestamp 1738175533
transform 1 0 27876 0 1 33184
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_57_290
timestamp 1738175533
transform 1 0 27784 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_314
timestamp 1738175533
transform 1 0 29992 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_326
timestamp 1738175533
transform 1 0 31096 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1738175533
transform 1 0 32568 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1738175533
transform 1 0 33396 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_338
timestamp 1738175533
transform 1 0 32200 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_343
timestamp 1738175533
transform 1 0 32660 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_354
timestamp 1738175533
transform 1 0 33672 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1738175533
transform -1 0 34316 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1738175533
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1738175533
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1738175533
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1738175533
transform 1 0 3772 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_27
timestamp 1738175533
transform 1 0 3588 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_30
timestamp 1738175533
transform 1 0 3864 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_42
timestamp 1738175533
transform 1 0 4968 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_54
timestamp 1738175533
transform 1 0 6072 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_66
timestamp 1738175533
transform 1 0 7176 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1642_
timestamp 1738175533
transform 1 0 9844 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1738175533
transform 1 0 9016 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_78
timestamp 1738175533
transform 1 0 8280 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_87
timestamp 1738175533
transform 1 0 9108 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_111
timestamp 1738175533
transform 1 0 11316 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_119
timestamp 1738175533
transform 1 0 12052 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1458_
timestamp 1738175533
transform 1 0 13432 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1569_
timestamp 1738175533
transform 1 0 12236 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1738175533
transform 1 0 14260 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_130
timestamp 1738175533
transform 1 0 13064 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_137
timestamp 1738175533
transform 1 0 13708 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_144
timestamp 1738175533
transform 1 0 14352 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_156
timestamp 1738175533
transform 1 0 15456 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__dfstp_1  _1745_
timestamp 1738175533
transform 1 0 17112 0 -1 34272
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_58_168
timestamp 1738175533
transform 1 0 16560 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1738175533
transform 1 0 19504 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_195
timestamp 1738175533
transform 1 0 19044 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_199
timestamp 1738175533
transform 1 0 19412 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_201
timestamp 1738175533
transform 1 0 19596 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_213
timestamp 1738175533
transform 1 0 20700 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _1748_
timestamp 1738175533
transform 1 0 20976 0 -1 34272
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_58_237
timestamp 1738175533
transform 1 0 22908 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1044_
timestamp 1738175533
transform 1 0 23276 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1738175533
transform 1 0 24748 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_250
timestamp 1738175533
transform 1 0 24104 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_256
timestamp 1738175533
transform 1 0 24656 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_258
timestamp 1738175533
transform 1 0 24840 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_270
timestamp 1738175533
transform 1 0 25944 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_282
timestamp 1738175533
transform 1 0 27048 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_294
timestamp 1738175533
transform 1 0 28152 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_306
timestamp 1738175533
transform 1 0 29256 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1738175533
transform 1 0 29992 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_315
timestamp 1738175533
transform 1 0 30084 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_327
timestamp 1738175533
transform 1 0 31188 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_339
timestamp 1738175533
transform 1 0 32292 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_351
timestamp 1738175533
transform 1 0 33396 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_357
timestamp 1738175533
transform 1 0 33948 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1738175533
transform -1 0 34316 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1738175533
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1738175533
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1738175533
transform -1 0 3036 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1738175533
transform 1 0 1380 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1738175533
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1738175533
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_7
timestamp 1738175533
transform 1 0 1748 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_15
timestamp 1738175533
transform 1 0 2484 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_21
timestamp 1738175533
transform 1 0 3036 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1738175533
transform 1 0 3772 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1738175533
transform -1 0 5336 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1738175533
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1738175533
transform 1 0 4692 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_30
timestamp 1738175533
transform 1 0 3864 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_42
timestamp 1738175533
transform 1 0 4968 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_46
timestamp 1738175533
transform 1 0 5336 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1583_
timestamp 1738175533
transform -1 0 8464 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1738175533
transform 1 0 6348 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1738175533
transform 1 0 6440 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1738175533
transform -1 0 7452 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_51
timestamp 1738175533
transform 1 0 5796 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_58
timestamp 1738175533
transform 1 0 6440 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_70
timestamp 1738175533
transform 1 0 7544 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_59
timestamp 1738175533
transform 1 0 6532 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_69
timestamp 1738175533
transform 1 0 7452 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1298_
timestamp 1738175533
transform 1 0 9660 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1584_
timestamp 1738175533
transform -1 0 8648 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1738175533
transform 1 0 9108 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_80
timestamp 1738175533
transform 1 0 8464 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_92
timestamp 1738175533
transform 1 0 9568 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_82
timestamp 1738175533
transform 1 0 8648 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_86
timestamp 1738175533
transform 1 0 9016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_88
timestamp 1738175533
transform 1 0 9200 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output24
timestamp 1738175533
transform -1 0 10948 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_100
timestamp 1738175533
transform 1 0 10304 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_107
timestamp 1738175533
transform 1 0 10948 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1570_
timestamp 1738175533
transform 1 0 12052 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1738175533
transform 1 0 11592 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1738175533
transform 1 0 11776 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_111
timestamp 1738175533
transform 1 0 11316 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_115
timestamp 1738175533
transform 1 0 11684 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_115
timestamp 1738175533
transform 1 0 11684 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_99
timestamp 1738175533
transform 1 0 10212 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_117
timestamp 1738175533
transform 1 0 11868 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1606_
timestamp 1738175533
transform 1 0 13800 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output23
timestamp 1738175533
transform -1 0 13708 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_128
timestamp 1738175533
transform 1 0 12880 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_136
timestamp 1738175533
transform 1 0 13616 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_129
timestamp 1738175533
transform 1 0 12972 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_137
timestamp 1738175533
transform 1 0 13708 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1738175533
transform 1 0 14444 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1738175533
transform 1 0 16100 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_154
timestamp 1738175533
transform 1 0 15272 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_166
timestamp 1738175533
transform 1 0 16376 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_146
timestamp 1738175533
transform 1 0 14536 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_158
timestamp 1738175533
transform 1 0 15640 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_162
timestamp 1738175533
transform 1 0 16008 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_166
timestamp 1738175533
transform 1 0 16376 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1738175533
transform 1 0 16836 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1738175533
transform 1 0 17112 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_170
timestamp 1738175533
transform 1 0 16744 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_172
timestamp 1738175533
transform 1 0 16928 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_184
timestamp 1738175533
transform 1 0 18032 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_175
timestamp 1738175533
transform 1 0 17204 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_187
timestamp 1738175533
transform 1 0 18308 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__dfstp_1  _1746_
timestamp 1738175533
transform 1 0 19044 0 1 34272
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1738175533
transform 1 0 19780 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1738175533
transform 1 0 18860 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_192
timestamp 1738175533
transform 1 0 18768 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_197
timestamp 1738175533
transform 1 0 19228 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_204
timestamp 1738175533
transform 1 0 19872 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output38
timestamp 1738175533
transform -1 0 21988 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_216
timestamp 1738175533
transform 1 0 20976 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_222
timestamp 1738175533
transform 1 0 21528 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1738175533
transform 1 0 22080 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1738175533
transform 1 0 22448 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_229
timestamp 1738175533
transform 1 0 22172 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_233
timestamp 1738175533
transform 1 0 22540 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_227
timestamp 1738175533
transform 1 0 21988 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_231
timestamp 1738175533
transform 1 0 22356 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _1749_
timestamp 1738175533
transform 1 0 22632 0 1 34272
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_59_216
timestamp 1738175533
transform 1 0 20976 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1738175533
transform 1 0 22540 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1738175533
transform 1 0 25116 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output25
timestamp 1738175533
transform -1 0 24748 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_255
timestamp 1738175533
transform 1 0 24564 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_245
timestamp 1738175533
transform 1 0 23644 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_257
timestamp 1738175533
transform 1 0 24748 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_262
timestamp 1738175533
transform 1 0 25208 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1738175533
transform 1 0 27324 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  input13
timestamp 1738175533
transform -1 0 27416 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_267
timestamp 1738175533
transform 1 0 25668 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_279
timestamp 1738175533
transform 1 0 26772 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_286
timestamp 1738175533
transform 1 0 27416 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_274
timestamp 1738175533
transform 1 0 26312 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_286
timestamp 1738175533
transform 1 0 27416 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1460_
timestamp 1738175533
transform -1 0 29532 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1738175533
transform 1 0 27784 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_298
timestamp 1738175533
transform 1 0 28520 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_309
timestamp 1738175533
transform 1 0 29532 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_291
timestamp 1738175533
transform 1 0 27876 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_303
timestamp 1738175533
transform 1 0 28980 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1738175533
transform 1 0 30452 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1738175533
transform 1 0 29808 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1738175533
transform -1 0 32016 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_321
timestamp 1738175533
transform 1 0 30636 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_333
timestamp 1738175533
transform 1 0 31740 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_311
timestamp 1738175533
transform 1 0 29716 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_315
timestamp 1738175533
transform 1 0 30084 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_320
timestamp 1738175533
transform 1 0 30544 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1738175533
transform 1 0 32568 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1738175533
transform -1 0 32752 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_341
timestamp 1738175533
transform 1 0 32476 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_336
timestamp 1738175533
transform 1 0 32016 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_344
timestamp 1738175533
transform 1 0 32752 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1738175533
transform 1 0 33120 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_355
timestamp 1738175533
transform 1 0 33764 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_349
timestamp 1738175533
transform 1 0 33212 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_357
timestamp 1738175533
transform 1 0 33948 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_343
timestamp 1738175533
transform 1 0 32660 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1738175533
transform -1 0 34316 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1738175533
transform -1 0 34316 0 -1 35360
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 16328 800 16448 4 clk_48
port 1 nsew
rlabel metal2 s 29918 36853 29974 37653 4 data_in[0]
port 2 nsew
rlabel metal3 s 0 8168 800 8288 4 data_in[1]
port 3 nsew
rlabel metal2 s 16118 36853 16174 37653 4 data_in[2]
port 4 nsew
rlabel metal2 s 13818 0 13874 800 4 data_in[3]
port 5 nsew
rlabel metal2 s 2778 36853 2834 37653 4 data_in[4]
port 6 nsew
rlabel metal3 s 34709 33328 35509 33448 4 data_in[5]
port 7 nsew
rlabel metal3 s 0 28568 800 28688 4 data_in[6]
port 8 nsew
rlabel metal3 s 34709 21088 35509 21208 4 data_in[7]
port 9 nsew
rlabel metal3 s 34709 25168 35509 25288 4 data_in_valid
port 10 nsew
rlabel metal2 s 13358 36853 13414 37653 4 data_out[0]
port 11 nsew
rlabel metal2 s 10598 36853 10654 37653 4 data_out[1]
port 12 nsew
rlabel metal2 s 24398 36853 24454 37653 4 data_out[2]
port 13 nsew
rlabel metal2 s 8298 0 8354 800 4 data_out[3]
port 14 nsew
rlabel metal2 s 27618 0 27674 800 4 data_out[4]
port 15 nsew
rlabel metal3 s 0 20408 800 20528 4 data_out[5]
port 16 nsew
rlabel metal2 s 19338 0 19394 800 4 data_out[6]
port 17 nsew
rlabel metal2 s 22098 0 22154 800 4 data_out[7]
port 18 nsew
rlabel metal3 s 0 4088 800 4208 4 data_strobe
port 19 nsew
rlabel metal2 s 7838 36853 7894 37653 4 data_toggle
port 20 nsew
rlabel metal2 s 478 0 534 800 4 direction_in
port 21 nsew
rlabel metal2 s 30378 0 30434 800 4 endpoint[0]
port 22 nsew
rlabel metal3 s 34709 12928 35509 13048 4 endpoint[1]
port 23 nsew
rlabel metal2 s 32678 0 32734 800 4 endpoint[2]
port 24 nsew
rlabel metal2 s 16578 0 16634 800 4 endpoint[3]
port 25 nsew
rlabel metal3 s 0 24488 800 24608 4 handshake[0]
port 26 nsew
rlabel metal3 s 0 32648 800 32768 4 handshake[1]
port 27 nsew
rlabel metal2 s 27158 36853 27214 37653 4 rst_n
port 28 nsew
rlabel metal2 s 5078 36853 5134 37653 4 rx_j
port 29 nsew
rlabel metal3 s 34709 29248 35509 29368 4 rx_se0
port 30 nsew
rlabel metal3 s 34709 688 35509 808 4 setup
port 31 nsew
rlabel metal2 s 21638 36853 21694 37653 4 success
port 32 nsew
rlabel metal2 s 11058 0 11114 800 4 transaction_active
port 33 nsew
rlabel metal3 s 34709 17008 35509 17128 4 tx_en
port 34 nsew
rlabel metal2 s 24858 0 24914 800 4 tx_j
port 35 nsew
rlabel metal3 s 0 12248 800 12368 4 tx_se0
port 36 nsew
rlabel metal2 s 5538 0 5594 800 4 usb_address[0]
port 37 nsew
rlabel metal2 s 32678 36853 32734 37653 4 usb_address[1]
port 38 nsew
rlabel metal2 s 18878 36853 18934 37653 4 usb_address[2]
port 39 nsew
rlabel metal3 s 34709 8848 35509 8968 4 usb_address[3]
port 40 nsew
rlabel metal3 s 0 36728 800 36848 4 usb_address[4]
port 41 nsew
rlabel metal2 s 2778 0 2834 800 4 usb_address[5]
port 42 nsew
rlabel metal2 s 34978 36853 35034 37653 4 usb_address[6]
port 43 nsew
rlabel metal3 s 34709 4768 35509 4888 4 usb_rst
port 44 nsew
rlabel metal4 s 28621 2128 28941 35408 4 VPWR
port 45 nsew
rlabel metal4 s 17550 2128 17870 35408 4 VPWR
port 45 nsew
rlabel metal4 s 6479 2128 6799 35408 4 VPWR
port 45 nsew
rlabel metal5 s 1104 29621 34316 29941 4 VPWR
port 45 nsew
rlabel metal5 s 1104 18560 34316 18880 4 VPWR
port 45 nsew
rlabel metal5 s 1104 7499 34316 7819 4 VPWR
port 45 nsew
rlabel metal4 s 23085 2128 23405 35408 4 VGND
port 46 nsew
rlabel metal4 s 12015 2128 12335 35408 4 VGND
port 46 nsew
rlabel metal5 s 1104 24091 34316 24411 4 VGND
port 46 nsew
rlabel metal5 s 1104 13029 34316 13349 4 VGND
port 46 nsew
<< properties >>
string FIXED_BBOX 0 0 35509 37653
<< end >>
